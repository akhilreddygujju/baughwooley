magic
tech scmos
timestamp 1733271326
<< polysilicon >>
rect 163 133 165 147
rect 18 81 20 100
rect 26 81 28 100
rect 64 87 66 99
rect 82 87 84 106
rect 100 87 102 99
rect 108 87 110 89
rect 116 87 118 99
rect 124 87 126 89
rect 145 87 147 129
rect 163 87 165 129
rect 181 87 183 99
rect 189 87 191 89
rect 197 87 199 99
rect 205 87 207 89
rect 227 87 229 107
rect 235 87 237 107
rect 251 87 253 89
rect 278 87 280 129
rect 286 87 288 147
rect 302 87 304 89
rect 324 87 326 99
rect 332 87 334 89
rect 355 87 357 89
rect 18 47 20 73
rect 26 47 28 73
rect 18 37 20 39
rect 26 37 28 39
rect 64 37 66 79
rect 82 37 84 79
rect 100 41 102 71
rect 108 41 110 71
rect 116 41 118 71
rect 124 41 126 71
rect 145 37 147 79
rect 163 37 165 79
rect 181 41 183 71
rect 189 41 191 71
rect 197 41 199 71
rect 205 41 207 71
rect 227 41 229 79
rect 235 41 237 79
rect 251 37 253 79
rect 278 41 280 79
rect 286 41 288 79
rect 302 37 304 79
rect 324 41 326 79
rect 332 41 334 79
rect 355 37 357 79
rect 64 31 66 33
rect 82 4 84 33
rect 100 31 102 33
rect 108 4 110 33
rect 116 31 118 33
rect 124 15 126 33
rect 145 31 147 33
rect 163 17 165 33
rect 181 31 183 33
rect 189 17 191 33
rect 197 31 199 33
rect 205 21 207 33
rect 227 31 229 33
rect 235 31 237 33
rect 251 31 253 33
rect 278 31 280 33
rect 286 31 288 33
rect 302 31 304 33
rect 324 31 326 33
rect 332 7 334 33
rect 355 31 357 33
<< ndiffusion >>
rect 17 39 18 47
rect 20 39 26 47
rect 28 39 29 47
rect 63 33 64 37
rect 66 33 67 37
rect 81 33 82 37
rect 84 33 85 37
rect 99 33 100 41
rect 102 33 108 41
rect 110 33 111 41
rect 115 33 116 41
rect 118 33 124 41
rect 126 33 127 41
rect 144 33 145 37
rect 147 33 148 37
rect 162 33 163 37
rect 165 33 166 37
rect 180 33 181 41
rect 183 33 189 41
rect 191 33 192 41
rect 196 33 197 41
rect 199 33 205 41
rect 207 33 208 41
rect 226 33 227 41
rect 229 33 235 41
rect 237 33 238 41
rect 250 33 251 37
rect 253 33 254 37
rect 277 33 278 41
rect 280 33 286 41
rect 288 33 289 41
rect 301 33 302 37
rect 304 33 305 37
rect 323 33 324 41
rect 326 33 327 41
rect 331 33 332 41
rect 334 33 335 41
rect 354 33 355 37
rect 357 33 358 37
<< pdiffusion >>
rect 17 73 18 81
rect 20 73 21 81
rect 25 73 26 81
rect 28 73 29 81
rect 63 79 64 87
rect 66 79 67 87
rect 81 79 82 87
rect 84 79 85 87
rect 99 71 100 87
rect 102 79 103 87
rect 107 79 108 87
rect 102 71 108 79
rect 110 71 111 87
rect 115 71 116 87
rect 118 79 124 87
rect 118 71 119 79
rect 123 71 124 79
rect 126 71 127 87
rect 144 79 145 87
rect 147 79 148 87
rect 162 79 163 87
rect 165 79 166 87
rect 180 71 181 87
rect 183 79 184 87
rect 188 79 189 87
rect 183 71 189 79
rect 191 71 192 87
rect 196 71 197 87
rect 199 79 205 87
rect 199 71 200 79
rect 204 71 205 79
rect 207 71 208 87
rect 226 79 227 87
rect 229 79 230 87
rect 234 79 235 87
rect 237 79 238 87
rect 250 79 251 87
rect 253 79 254 87
rect 277 79 278 87
rect 280 79 281 87
rect 285 79 286 87
rect 288 79 289 87
rect 301 79 302 87
rect 304 79 305 87
rect 323 79 324 87
rect 326 79 332 87
rect 334 79 335 87
rect 354 79 355 87
rect 357 79 358 87
<< metal1 >>
rect 166 147 285 151
rect 63 122 230 126
rect 63 103 67 122
rect 81 110 85 113
rect 226 111 230 122
rect 234 111 238 114
rect 67 99 99 103
rect 112 99 115 103
rect 151 99 180 103
rect 193 99 196 103
rect 316 99 323 103
rect 13 95 362 96
rect 13 91 21 95
rect 25 91 73 95
rect 77 91 156 95
rect 160 91 230 95
rect 234 91 247 95
rect 251 91 281 95
rect 285 91 298 95
rect 302 91 327 95
rect 331 91 351 95
rect 355 91 362 95
rect 13 90 362 91
rect 13 81 17 90
rect 29 81 33 90
rect 59 87 63 90
rect 77 87 81 90
rect 103 87 107 90
rect 140 87 144 90
rect 158 87 162 90
rect 184 87 188 90
rect 222 87 226 90
rect 238 87 242 90
rect 21 62 25 73
rect 67 64 71 79
rect 85 64 89 79
rect 99 71 111 75
rect 115 83 127 87
rect 21 61 33 62
rect 21 58 60 61
rect 29 57 60 58
rect 119 59 123 71
rect 148 64 152 79
rect 166 64 170 79
rect 180 71 192 75
rect 196 83 208 87
rect 246 87 250 90
rect 273 87 277 90
rect 289 87 293 90
rect 297 87 301 90
rect 319 87 323 90
rect 350 87 354 90
rect 200 59 204 71
rect 230 64 234 79
rect 254 64 258 79
rect 281 64 285 79
rect 305 64 309 79
rect 335 64 339 79
rect 230 60 247 64
rect 29 47 33 57
rect 13 30 17 39
rect 67 37 71 59
rect 85 37 89 59
rect 111 55 141 59
rect 111 41 115 55
rect 148 37 152 59
rect 166 37 170 59
rect 192 55 214 59
rect 192 41 196 55
rect 238 41 242 60
rect 59 30 63 33
rect 77 30 81 33
rect 95 30 99 33
rect 127 30 131 33
rect 140 30 144 33
rect 158 30 162 33
rect 176 30 180 33
rect 208 30 212 33
rect 281 60 298 64
rect 254 37 258 59
rect 289 41 293 60
rect 327 60 351 64
rect 305 37 309 59
rect 327 41 331 60
rect 358 37 362 79
rect 222 30 226 33
rect 246 30 250 33
rect 273 30 277 33
rect 297 30 301 33
rect 319 30 323 33
rect 335 30 339 33
rect 350 30 354 33
rect 13 29 362 30
rect 13 25 14 29
rect 18 25 60 29
rect 64 25 141 29
rect 145 25 223 29
rect 227 25 247 29
rect 251 25 274 29
rect 278 25 298 29
rect 302 25 320 29
rect 324 25 351 29
rect 355 25 362 29
rect 13 24 362 25
rect 120 11 123 15
rect 166 13 188 17
rect 201 17 204 21
rect 85 0 107 4
rect 327 3 331 7
<< metal2 >>
rect 148 129 277 133
rect 86 114 234 118
rect 107 96 111 99
rect 188 96 192 99
rect 311 96 315 99
rect 86 92 111 96
rect 167 92 192 96
rect 255 92 315 96
rect 86 64 90 92
rect 167 64 171 92
rect 255 64 259 92
rect 68 28 72 59
rect 149 28 153 59
rect 68 24 119 28
rect 149 24 200 28
rect 115 15 119 24
rect 196 21 200 24
rect 306 7 310 59
rect 306 3 322 7
<< ntransistor >>
rect 18 39 20 47
rect 26 39 28 47
rect 64 33 66 37
rect 82 33 84 37
rect 100 33 102 41
rect 108 33 110 41
rect 116 33 118 41
rect 124 33 126 41
rect 145 33 147 37
rect 163 33 165 37
rect 181 33 183 41
rect 189 33 191 41
rect 197 33 199 41
rect 205 33 207 41
rect 227 33 229 41
rect 235 33 237 41
rect 251 33 253 37
rect 278 33 280 41
rect 286 33 288 41
rect 302 33 304 37
rect 324 33 326 41
rect 332 33 334 41
rect 355 33 357 37
<< ptransistor >>
rect 18 73 20 81
rect 26 73 28 81
rect 64 79 66 87
rect 82 79 84 87
rect 100 71 102 87
rect 108 71 110 87
rect 116 71 118 87
rect 124 71 126 87
rect 145 79 147 87
rect 163 79 165 87
rect 181 71 183 87
rect 189 71 191 87
rect 197 71 199 87
rect 205 71 207 87
rect 227 79 229 87
rect 235 79 237 87
rect 251 79 253 87
rect 278 79 280 87
rect 286 79 288 87
rect 302 79 304 87
rect 324 79 326 87
rect 332 79 334 87
rect 355 79 357 87
<< polycontact >>
rect 162 147 166 151
rect 285 147 289 151
rect 144 129 148 133
rect 277 129 281 133
rect 81 106 85 110
rect 17 100 21 104
rect 25 100 29 104
rect 63 99 67 103
rect 99 99 103 103
rect 115 99 119 103
rect 147 99 151 103
rect 226 107 230 111
rect 234 107 238 111
rect 180 99 184 103
rect 196 99 200 103
rect 323 99 327 103
rect 60 57 64 61
rect 78 60 82 64
rect 141 55 145 59
rect 247 60 251 64
rect 298 60 302 64
rect 351 60 355 64
rect 204 17 208 21
rect 123 11 127 15
rect 162 13 166 17
rect 188 13 192 17
rect 81 0 85 4
rect 107 0 111 4
rect 331 3 335 7
<< ndcontact >>
rect 13 39 17 47
rect 29 39 33 47
rect 59 33 63 37
rect 67 33 71 37
rect 77 33 81 37
rect 85 33 89 37
rect 95 33 99 41
rect 111 33 115 41
rect 127 33 131 41
rect 140 33 144 37
rect 148 33 152 37
rect 158 33 162 37
rect 166 33 170 37
rect 176 33 180 41
rect 192 33 196 41
rect 208 33 212 41
rect 222 33 226 41
rect 238 33 242 41
rect 246 33 250 37
rect 254 33 258 37
rect 273 33 277 41
rect 289 33 293 41
rect 297 33 301 37
rect 305 33 309 37
rect 319 33 323 41
rect 327 33 331 41
rect 335 33 339 41
rect 350 33 354 37
rect 358 33 362 37
<< pdcontact >>
rect 13 73 17 81
rect 21 73 25 81
rect 29 73 33 81
rect 59 79 63 87
rect 67 79 71 87
rect 77 79 81 87
rect 85 79 89 87
rect 95 71 99 87
rect 103 79 107 87
rect 111 71 115 87
rect 119 71 123 79
rect 127 71 131 87
rect 140 79 144 87
rect 148 79 152 87
rect 158 79 162 87
rect 166 79 170 87
rect 176 71 180 87
rect 184 79 188 87
rect 192 71 196 87
rect 200 71 204 79
rect 208 71 212 87
rect 222 79 226 87
rect 230 79 234 87
rect 238 79 242 87
rect 246 79 250 87
rect 254 79 258 87
rect 273 79 277 87
rect 281 79 285 87
rect 289 79 293 87
rect 297 79 301 87
rect 305 79 309 87
rect 319 79 323 87
rect 335 79 339 87
rect 350 79 354 87
rect 358 79 362 87
<< m2contact >>
rect 81 113 86 118
rect 234 114 239 119
rect 107 99 112 104
rect 188 99 193 104
rect 311 99 316 104
rect 67 59 72 64
rect 85 59 90 64
rect 148 59 153 64
rect 166 59 171 64
rect 254 59 259 64
rect 305 59 310 64
rect 115 10 120 15
rect 196 16 201 21
rect 322 2 327 7
<< psubstratepcontact >>
rect 14 25 18 29
rect 60 25 64 29
rect 141 25 145 29
rect 223 25 227 29
rect 247 25 251 29
rect 274 25 278 29
rect 298 25 302 29
rect 320 25 324 29
rect 351 25 355 29
<< nsubstratencontact >>
rect 21 91 25 95
rect 73 91 77 95
rect 156 91 160 95
rect 230 91 234 95
rect 247 91 251 95
rect 281 91 285 95
rect 298 91 302 95
rect 327 91 331 95
rect 351 91 355 95
<< labels >>
rlabel metal1 174 93 174 93 5 vdd
rlabel metal1 174 27 174 27 1 gnd
rlabel metal1 211 57 211 57 1 S
rlabel polycontact 80 62 80 62 1 B
rlabel m2contact 69 61 69 61 1 not1_1
rlabel m2contact 87 61 87 61 1 not1_2
rlabel m2contact 150 62 150 62 1 not2_1
rlabel m2contact 168 61 168 61 1 not2_2
rlabel polycontact 143 57 143 57 1 out_XOR1
rlabel polycontact 249 62 249 62 1 out_AND1
rlabel polycontact 300 62 300 62 1 out_AND2
rlabel polycontact 353 62 353 62 1 out_OR
rlabel metal1 360 62 360 62 7 cout
rlabel polycontact 164 149 164 149 5 cin
rlabel polycontact 19 102 19 102 1 X
rlabel polycontact 27 102 27 102 1 Y
rlabel polycontact 62 59 62 59 1 A
<< end >>
