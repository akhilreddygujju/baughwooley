magic
tech scmos
timestamp 1733699845
<< polysilicon >>
rect -54 81 -52 110
rect -46 81 -44 110
rect 2 97 4 110
rect 18 97 20 99
rect 34 97 36 110
rect 42 97 44 99
rect 50 97 52 110
rect 58 97 60 99
rect 77 97 79 109
rect 85 97 87 109
rect 103 97 105 99
rect 131 97 133 110
rect 147 97 149 99
rect 163 97 165 110
rect 171 97 173 99
rect 179 97 181 110
rect 187 97 189 99
rect 206 97 208 109
rect 214 97 216 109
rect 232 97 234 99
rect 259 97 261 109
rect 267 97 269 109
rect 285 97 287 99
rect -30 81 -28 83
rect -54 47 -52 73
rect -46 47 -44 73
rect -30 43 -28 73
rect -54 37 -52 39
rect -46 37 -44 39
rect -30 37 -28 39
rect 2 29 4 89
rect 18 29 20 89
rect 34 33 36 81
rect 42 33 44 81
rect 50 33 52 81
rect 58 33 60 81
rect 77 33 79 89
rect 85 33 87 89
rect 103 29 105 89
rect 131 29 133 89
rect 147 29 149 89
rect 163 33 165 81
rect 171 33 173 81
rect 179 33 181 81
rect 187 33 189 81
rect 206 33 208 89
rect 214 33 216 89
rect 232 29 234 89
rect 259 34 261 89
rect 267 34 269 89
rect 285 29 287 89
rect 2 23 4 25
rect 18 12 20 25
rect 34 23 36 25
rect 42 12 44 25
rect 50 23 52 25
rect 58 12 60 25
rect 77 23 79 25
rect 85 13 87 25
rect 103 23 105 25
rect 131 23 133 25
rect 147 12 149 25
rect 163 23 165 25
rect 171 12 173 25
rect 179 23 181 25
rect 187 12 189 25
rect 206 23 208 25
rect 214 13 216 25
rect 232 23 234 25
rect 259 23 261 26
rect 267 13 269 26
rect 285 23 287 25
<< ndiffusion >>
rect -55 39 -54 47
rect -52 39 -46 47
rect -44 39 -43 47
rect -31 39 -30 43
rect -28 39 -27 43
rect 1 25 2 29
rect 4 25 5 29
rect 17 25 18 29
rect 20 25 21 29
rect 33 25 34 33
rect 36 25 42 33
rect 44 25 45 33
rect 49 25 50 33
rect 52 25 58 33
rect 60 25 61 33
rect 74 25 77 33
rect 79 25 85 33
rect 87 25 90 33
rect 102 25 103 29
rect 105 25 106 29
rect 130 25 131 29
rect 133 25 134 29
rect 146 25 147 29
rect 149 25 150 29
rect 162 25 163 33
rect 165 25 171 33
rect 173 25 174 33
rect 178 25 179 33
rect 181 25 187 33
rect 189 25 190 33
rect 203 25 206 33
rect 208 25 214 33
rect 216 25 219 33
rect 231 25 232 29
rect 234 25 235 29
rect 257 26 259 34
rect 261 26 262 34
rect 266 26 267 34
rect 269 26 270 34
rect 283 25 285 29
rect 287 25 289 29
<< pdiffusion >>
rect 1 89 2 97
rect 4 89 5 97
rect 17 89 18 97
rect 20 89 21 97
rect -55 73 -54 81
rect -52 73 -51 81
rect -47 73 -46 81
rect -44 73 -43 81
rect -31 73 -30 81
rect -28 73 -27 81
rect 33 81 34 97
rect 36 89 37 97
rect 41 89 42 97
rect 36 81 42 89
rect 44 81 45 97
rect 49 81 50 97
rect 52 89 58 97
rect 52 81 53 89
rect 57 81 58 89
rect 60 81 61 97
rect 70 95 77 97
rect 70 91 71 95
rect 75 91 77 95
rect 70 89 77 91
rect 79 95 85 97
rect 79 91 80 95
rect 84 91 85 95
rect 79 89 85 91
rect 87 95 94 97
rect 87 91 89 95
rect 93 91 94 95
rect 87 89 94 91
rect 102 89 103 97
rect 105 89 106 97
rect 130 89 131 97
rect 133 89 134 97
rect 146 89 147 97
rect 149 89 150 97
rect 162 81 163 97
rect 165 89 166 97
rect 170 89 171 97
rect 165 81 171 89
rect 173 81 174 97
rect 178 81 179 97
rect 181 89 187 97
rect 181 81 182 89
rect 186 81 187 89
rect 189 81 190 97
rect 199 95 206 97
rect 199 91 200 95
rect 204 91 206 95
rect 199 89 206 91
rect 208 95 214 97
rect 208 91 209 95
rect 213 91 214 95
rect 208 89 214 91
rect 216 95 223 97
rect 216 91 218 95
rect 222 91 223 95
rect 216 89 223 91
rect 231 89 232 97
rect 234 89 235 97
rect 257 89 259 97
rect 261 89 267 97
rect 269 89 270 97
rect 283 89 285 97
rect 287 89 289 97
<< metal1 >>
rect 33 120 80 124
rect 33 114 37 120
rect 5 110 33 114
rect 46 110 49 114
rect 76 113 80 120
rect 162 120 209 124
rect 162 114 166 120
rect 134 110 162 114
rect 175 110 178 114
rect 205 113 209 120
rect -59 105 293 106
rect -59 101 -51 105
rect -47 101 -34 105
rect -30 101 14 105
rect 18 101 72 105
rect 76 101 89 105
rect 93 101 143 105
rect 147 101 201 105
rect 205 101 218 105
rect 222 101 254 105
rect 258 101 279 105
rect 283 101 293 105
rect -59 100 293 101
rect -59 81 -55 100
rect -43 81 -39 100
rect -35 81 -31 100
rect -3 97 1 100
rect 13 97 17 100
rect 37 97 41 100
rect -51 62 -47 73
rect -51 59 -39 62
rect -27 61 -23 73
rect 5 61 9 89
rect 21 61 25 89
rect 33 81 45 85
rect 49 93 61 97
rect 71 95 75 100
rect 89 95 93 100
rect 98 97 102 100
rect 126 97 130 100
rect 142 97 146 100
rect 166 97 170 100
rect 53 67 57 81
rect 45 63 65 67
rect -51 58 -34 59
rect -43 55 -34 58
rect -27 57 -2 61
rect -43 47 -39 55
rect -27 43 -23 57
rect -59 22 -55 39
rect -35 22 -31 39
rect 5 29 9 56
rect 21 29 25 56
rect 45 33 49 63
rect 80 58 84 91
rect 106 58 110 89
rect 125 77 127 81
rect 134 61 138 89
rect 150 61 154 89
rect 162 81 174 85
rect 178 93 190 97
rect 200 95 204 100
rect 218 95 222 100
rect 227 97 231 100
rect 253 97 257 100
rect 279 97 283 100
rect 182 67 186 81
rect 174 63 194 67
rect 80 54 99 58
rect 106 54 113 58
rect 90 33 94 54
rect -3 22 1 25
rect 13 22 17 25
rect 29 22 33 25
rect 61 22 65 25
rect 106 29 110 54
rect 134 29 138 56
rect 150 29 154 56
rect 174 33 178 63
rect 209 58 213 91
rect 235 58 239 89
rect 270 84 274 89
rect 289 84 293 89
rect 262 80 281 84
rect 289 80 297 84
rect 209 54 228 58
rect 235 54 255 58
rect 219 33 223 54
rect 70 22 74 25
rect 98 22 102 25
rect 126 22 130 25
rect 142 22 146 25
rect 158 22 162 25
rect 190 22 194 25
rect 235 29 239 54
rect 262 34 266 80
rect 289 29 293 80
rect 199 22 203 25
rect 227 22 231 25
rect 253 22 257 26
rect 270 22 274 26
rect 279 22 283 25
rect -59 21 293 22
rect -59 17 -58 21
rect -54 17 -34 21
rect -30 17 -2 21
rect 2 17 71 21
rect 75 17 89 21
rect 93 17 99 21
rect 103 17 127 21
rect 131 17 200 21
rect 204 17 218 21
rect 222 17 228 21
rect 232 17 261 21
rect 265 17 279 21
rect 283 17 293 21
rect -59 16 293 17
rect 21 8 41 12
rect 41 1 45 8
rect 54 8 57 12
rect 84 1 88 9
rect 150 8 170 12
rect 41 -3 88 1
rect 170 1 174 8
rect 183 8 186 12
rect 213 1 217 9
rect 266 7 270 9
rect 170 -3 217 1
<< metal2 >>
rect 42 106 46 110
rect 171 106 175 110
rect 22 102 46 106
rect 151 102 175 106
rect 22 61 26 102
rect 120 66 124 76
rect 70 62 124 66
rect 151 61 155 102
rect 199 62 298 66
rect 6 20 10 56
rect 6 16 53 20
rect 49 12 53 16
rect 114 -5 118 53
rect 135 20 139 56
rect 135 16 182 20
rect 178 12 182 16
rect 265 -5 269 2
rect 114 -9 269 -5
<< ntransistor >>
rect -54 39 -52 47
rect -46 39 -44 47
rect -30 39 -28 43
rect 2 25 4 29
rect 18 25 20 29
rect 34 25 36 33
rect 42 25 44 33
rect 50 25 52 33
rect 58 25 60 33
rect 77 25 79 33
rect 85 25 87 33
rect 103 25 105 29
rect 131 25 133 29
rect 147 25 149 29
rect 163 25 165 33
rect 171 25 173 33
rect 179 25 181 33
rect 187 25 189 33
rect 206 25 208 33
rect 214 25 216 33
rect 232 25 234 29
rect 259 26 261 34
rect 267 26 269 34
rect 285 25 287 29
<< ptransistor >>
rect 2 89 4 97
rect 18 89 20 97
rect -54 73 -52 81
rect -46 73 -44 81
rect -30 73 -28 81
rect 34 81 36 97
rect 42 81 44 97
rect 50 81 52 97
rect 58 81 60 97
rect 77 89 79 97
rect 85 89 87 97
rect 103 89 105 97
rect 131 89 133 97
rect 147 89 149 97
rect 163 81 165 97
rect 171 81 173 97
rect 179 81 181 97
rect 187 81 189 97
rect 206 89 208 97
rect 214 89 216 97
rect 232 89 234 97
rect 259 89 261 97
rect 267 89 269 97
rect 285 89 287 97
<< polycontact >>
rect -55 110 -51 114
rect -47 110 -43 114
rect 1 110 5 114
rect 33 110 37 114
rect 49 110 53 114
rect 76 109 80 113
rect 130 110 134 114
rect 162 110 166 114
rect 178 110 182 114
rect 205 109 209 113
rect -34 55 -30 59
rect -2 57 2 61
rect 14 77 18 81
rect 99 54 103 58
rect 127 77 131 81
rect 143 77 147 81
rect 228 54 232 58
rect 255 54 259 58
rect 281 80 285 84
rect 17 8 21 12
rect 41 8 45 12
rect 57 8 61 12
rect 84 9 88 13
rect 146 8 150 12
rect 170 8 174 12
rect 186 8 190 12
rect 213 9 217 13
rect 266 9 270 13
<< ndcontact >>
rect -59 39 -55 47
rect -43 39 -39 47
rect -35 39 -31 43
rect -27 39 -23 43
rect -3 25 1 29
rect 5 25 9 29
rect 13 25 17 29
rect 21 25 25 29
rect 29 25 33 33
rect 45 25 49 33
rect 61 25 65 33
rect 70 25 74 33
rect 90 25 94 33
rect 98 25 102 29
rect 106 25 110 29
rect 126 25 130 29
rect 134 25 138 29
rect 142 25 146 29
rect 150 25 154 29
rect 158 25 162 33
rect 174 25 178 33
rect 190 25 194 33
rect 199 25 203 33
rect 219 25 223 33
rect 227 25 231 29
rect 235 25 239 29
rect 253 26 257 34
rect 262 26 266 34
rect 270 26 274 34
rect 279 25 283 29
rect 289 25 293 29
<< pdcontact >>
rect -3 89 1 97
rect 5 89 9 97
rect 13 89 17 97
rect 21 89 25 97
rect -59 73 -55 81
rect -51 73 -47 81
rect -43 73 -39 81
rect -35 73 -31 81
rect -27 73 -23 81
rect 29 81 33 97
rect 37 89 41 97
rect 45 81 49 97
rect 53 81 57 89
rect 61 81 65 97
rect 71 91 75 95
rect 80 91 84 95
rect 89 91 93 95
rect 98 89 102 97
rect 106 89 110 97
rect 126 89 130 97
rect 134 89 138 97
rect 142 89 146 97
rect 150 89 154 97
rect 158 81 162 97
rect 166 89 170 97
rect 174 81 178 97
rect 182 81 186 89
rect 190 81 194 97
rect 200 91 204 95
rect 209 91 213 95
rect 218 91 222 95
rect 227 89 231 97
rect 235 89 239 97
rect 253 89 257 97
rect 270 89 274 97
rect 279 89 283 97
rect 289 89 293 97
<< m2contact >>
rect 41 110 46 115
rect 170 110 175 115
rect 5 56 10 61
rect 21 56 26 61
rect 65 62 70 67
rect 120 76 125 81
rect 113 53 118 58
rect 134 56 139 61
rect 150 56 155 61
rect 194 62 199 67
rect 49 7 54 12
rect 178 7 183 12
rect 265 2 270 7
<< psubstratepcontact >>
rect -58 17 -54 21
rect -34 17 -30 21
rect -2 17 2 21
rect 71 17 75 21
rect 89 17 93 21
rect 99 17 103 21
rect 127 17 131 21
rect 200 17 204 21
rect 218 17 222 21
rect 228 17 232 21
rect 261 17 265 21
rect 279 17 283 21
<< nsubstratencontact >>
rect -51 101 -47 105
rect -34 101 -30 105
rect 14 101 18 105
rect 72 101 76 105
rect 89 101 93 105
rect 143 101 147 105
rect 201 101 205 105
rect 218 101 222 105
rect 254 101 258 105
rect 279 101 283 105
<< labels >>
rlabel metal1 -25 57 -25 57 7 vout
rlabel polycontact 16 79 16 79 1 B
rlabel polycontact 145 79 145 79 1 C
rlabel metal1 295 82 295 82 7 carry
rlabel metal2 296 64 296 64 7 sum
rlabel metal1 115 103 115 103 1 VDD
rlabel metal1 111 19 111 19 1 GND
rlabel polycontact 0 59 0 59 3 A
rlabel polycontact -45 112 -45 112 1 Y
rlabel polycontact -53 112 -53 112 1 X
<< end >>
