magic
tech scmos
timestamp 1700524122
<< polysilicon >>
rect 6 100 8 113
rect 22 100 24 102
rect 38 100 40 113
rect 46 100 48 102
rect 54 100 56 113
rect 62 100 64 102
rect 81 100 83 112
rect 89 100 91 112
rect 107 100 109 102
rect 135 100 137 113
rect 151 100 153 102
rect 167 100 169 113
rect 175 100 177 102
rect 183 100 185 113
rect 191 100 193 102
rect 210 100 212 112
rect 218 100 220 112
rect 236 100 238 102
rect 263 100 265 112
rect 271 100 273 112
rect 289 100 291 102
rect 6 32 8 92
rect 22 32 24 92
rect 38 36 40 84
rect 46 36 48 84
rect 54 36 56 84
rect 62 36 64 84
rect 81 36 83 92
rect 89 36 91 92
rect 107 32 109 92
rect 135 32 137 92
rect 151 32 153 92
rect 167 36 169 84
rect 175 36 177 84
rect 183 36 185 84
rect 191 36 193 84
rect 210 36 212 92
rect 218 36 220 92
rect 236 32 238 92
rect 263 37 265 92
rect 271 37 273 92
rect 289 32 291 92
rect 6 26 8 28
rect 22 15 24 28
rect 38 26 40 28
rect 46 15 48 28
rect 54 26 56 28
rect 62 15 64 28
rect 81 26 83 28
rect 89 16 91 28
rect 107 26 109 28
rect 135 26 137 28
rect 151 15 153 28
rect 167 26 169 28
rect 175 15 177 28
rect 183 26 185 28
rect 191 15 193 28
rect 210 26 212 28
rect 218 16 220 28
rect 236 26 238 28
rect 263 26 265 29
rect 271 16 273 29
rect 289 26 291 28
<< ndiffusion >>
rect 5 28 6 32
rect 8 28 9 32
rect 21 28 22 32
rect 24 28 25 32
rect 37 28 38 36
rect 40 28 46 36
rect 48 28 49 36
rect 53 28 54 36
rect 56 28 62 36
rect 64 28 65 36
rect 78 28 81 36
rect 83 28 89 36
rect 91 28 94 36
rect 106 28 107 32
rect 109 28 110 32
rect 134 28 135 32
rect 137 28 138 32
rect 150 28 151 32
rect 153 28 154 32
rect 166 28 167 36
rect 169 28 175 36
rect 177 28 178 36
rect 182 28 183 36
rect 185 28 191 36
rect 193 28 194 36
rect 207 28 210 36
rect 212 28 218 36
rect 220 28 223 36
rect 235 28 236 32
rect 238 28 239 32
rect 261 29 263 37
rect 265 29 266 37
rect 270 29 271 37
rect 273 29 274 37
rect 287 28 289 32
rect 291 28 293 32
<< pdiffusion >>
rect 5 92 6 100
rect 8 92 9 100
rect 21 92 22 100
rect 24 92 25 100
rect 37 84 38 100
rect 40 92 41 100
rect 45 92 46 100
rect 40 84 46 92
rect 48 84 49 100
rect 53 84 54 100
rect 56 92 62 100
rect 56 84 57 92
rect 61 84 62 92
rect 64 84 65 100
rect 74 98 81 100
rect 74 94 75 98
rect 79 94 81 98
rect 74 92 81 94
rect 83 98 89 100
rect 83 94 84 98
rect 88 94 89 98
rect 83 92 89 94
rect 91 98 98 100
rect 91 94 93 98
rect 97 94 98 98
rect 91 92 98 94
rect 106 92 107 100
rect 109 92 110 100
rect 134 92 135 100
rect 137 92 138 100
rect 150 92 151 100
rect 153 92 154 100
rect 166 84 167 100
rect 169 92 170 100
rect 174 92 175 100
rect 169 84 175 92
rect 177 84 178 100
rect 182 84 183 100
rect 185 92 191 100
rect 185 84 186 92
rect 190 84 191 92
rect 193 84 194 100
rect 203 98 210 100
rect 203 94 204 98
rect 208 94 210 98
rect 203 92 210 94
rect 212 98 218 100
rect 212 94 213 98
rect 217 94 218 98
rect 212 92 218 94
rect 220 98 227 100
rect 220 94 222 98
rect 226 94 227 98
rect 220 92 227 94
rect 235 92 236 100
rect 238 92 239 100
rect 261 92 263 100
rect 265 92 271 100
rect 273 92 274 100
rect 287 92 289 100
rect 291 92 293 100
<< metal1 >>
rect 37 123 84 127
rect 37 117 41 123
rect 9 113 37 117
rect 50 113 53 117
rect 80 116 84 123
rect 166 123 213 127
rect 166 117 170 123
rect 138 113 166 117
rect 179 113 182 117
rect 209 116 213 123
rect 1 108 297 109
rect 1 104 18 108
rect 22 104 76 108
rect 80 104 93 108
rect 97 104 147 108
rect 151 104 205 108
rect 209 104 222 108
rect 226 104 258 108
rect 262 104 283 108
rect 287 104 297 108
rect 1 103 297 104
rect 1 100 5 103
rect 17 100 21 103
rect 41 100 45 103
rect 9 64 13 92
rect 25 64 29 92
rect 37 84 49 88
rect 53 96 65 100
rect 75 98 79 103
rect 93 98 97 103
rect 102 100 106 103
rect 130 100 134 103
rect 146 100 150 103
rect 170 100 174 103
rect 57 70 61 84
rect 49 66 69 70
rect 9 32 13 59
rect 25 32 29 59
rect 49 36 53 66
rect 84 61 88 94
rect 110 61 114 92
rect 129 80 131 84
rect 138 64 142 92
rect 154 64 158 92
rect 166 84 178 88
rect 182 96 194 100
rect 204 98 208 103
rect 222 98 226 103
rect 231 100 235 103
rect 257 100 261 103
rect 283 100 287 103
rect 186 70 190 84
rect 178 66 198 70
rect 84 57 103 61
rect 110 57 117 61
rect 94 36 98 57
rect 1 25 5 28
rect 17 25 21 28
rect 33 25 37 28
rect 65 25 69 28
rect 110 32 114 57
rect 138 32 142 59
rect 154 32 158 59
rect 178 36 182 66
rect 213 61 217 94
rect 239 61 243 92
rect 274 87 278 92
rect 293 87 297 92
rect 266 83 285 87
rect 293 83 301 87
rect 213 57 232 61
rect 239 57 259 61
rect 223 36 227 57
rect 74 25 78 28
rect 102 25 106 28
rect 130 25 134 28
rect 146 25 150 28
rect 162 25 166 28
rect 194 25 198 28
rect 239 32 243 57
rect 266 37 270 83
rect 293 32 297 83
rect 203 25 207 28
rect 231 25 235 28
rect 257 25 261 29
rect 274 25 278 29
rect 283 25 287 28
rect 0 24 297 25
rect 0 20 2 24
rect 6 20 75 24
rect 79 20 93 24
rect 97 20 103 24
rect 107 20 131 24
rect 135 20 204 24
rect 208 20 222 24
rect 226 20 232 24
rect 236 20 265 24
rect 269 20 283 24
rect 287 20 297 24
rect 0 19 297 20
rect 25 11 45 15
rect 45 4 49 11
rect 58 11 61 15
rect 88 4 92 12
rect 154 11 174 15
rect 45 0 92 4
rect 174 4 178 11
rect 187 11 190 15
rect 217 4 221 12
rect 270 10 274 12
rect 174 0 221 4
<< metal2 >>
rect 46 109 50 113
rect 175 109 179 113
rect 26 105 50 109
rect 155 105 179 109
rect 26 64 30 105
rect 124 69 128 79
rect 74 65 128 69
rect 155 64 159 105
rect 203 65 302 69
rect 10 23 14 59
rect 10 19 57 23
rect 53 15 57 19
rect 118 -2 122 56
rect 139 23 143 59
rect 139 19 186 23
rect 182 15 186 19
rect 269 -2 273 5
rect 118 -6 273 -2
<< ntransistor >>
rect 6 28 8 32
rect 22 28 24 32
rect 38 28 40 36
rect 46 28 48 36
rect 54 28 56 36
rect 62 28 64 36
rect 81 28 83 36
rect 89 28 91 36
rect 107 28 109 32
rect 135 28 137 32
rect 151 28 153 32
rect 167 28 169 36
rect 175 28 177 36
rect 183 28 185 36
rect 191 28 193 36
rect 210 28 212 36
rect 218 28 220 36
rect 236 28 238 32
rect 263 29 265 37
rect 271 29 273 37
rect 289 28 291 32
<< ptransistor >>
rect 6 92 8 100
rect 22 92 24 100
rect 38 84 40 100
rect 46 84 48 100
rect 54 84 56 100
rect 62 84 64 100
rect 81 92 83 100
rect 89 92 91 100
rect 107 92 109 100
rect 135 92 137 100
rect 151 92 153 100
rect 167 84 169 100
rect 175 84 177 100
rect 183 84 185 100
rect 191 84 193 100
rect 210 92 212 100
rect 218 92 220 100
rect 236 92 238 100
rect 263 92 265 100
rect 271 92 273 100
rect 289 92 291 100
<< polycontact >>
rect 5 113 9 117
rect 37 113 41 117
rect 53 113 57 117
rect 80 112 84 116
rect 134 113 138 117
rect 166 113 170 117
rect 182 113 186 117
rect 209 112 213 116
rect 2 80 6 84
rect 18 80 22 84
rect 103 57 107 61
rect 131 80 135 84
rect 147 80 151 84
rect 232 57 236 61
rect 259 57 263 61
rect 285 83 289 87
rect 21 11 25 15
rect 45 11 49 15
rect 61 11 65 15
rect 88 12 92 16
rect 150 11 154 15
rect 174 11 178 15
rect 190 11 194 15
rect 217 12 221 16
rect 270 12 274 16
<< ndcontact >>
rect 1 28 5 32
rect 9 28 13 32
rect 17 28 21 32
rect 25 28 29 32
rect 33 28 37 36
rect 49 28 53 36
rect 65 28 69 36
rect 74 28 78 36
rect 94 28 98 36
rect 102 28 106 32
rect 110 28 114 32
rect 130 28 134 32
rect 138 28 142 32
rect 146 28 150 32
rect 154 28 158 32
rect 162 28 166 36
rect 178 28 182 36
rect 194 28 198 36
rect 203 28 207 36
rect 223 28 227 36
rect 231 28 235 32
rect 239 28 243 32
rect 257 29 261 37
rect 266 29 270 37
rect 274 29 278 37
rect 283 28 287 32
rect 293 28 297 32
<< pdcontact >>
rect 1 92 5 100
rect 9 92 13 100
rect 17 92 21 100
rect 25 92 29 100
rect 33 84 37 100
rect 41 92 45 100
rect 49 84 53 100
rect 57 84 61 92
rect 65 84 69 100
rect 75 94 79 98
rect 84 94 88 98
rect 93 94 97 98
rect 102 92 106 100
rect 110 92 114 100
rect 130 92 134 100
rect 138 92 142 100
rect 146 92 150 100
rect 154 92 158 100
rect 162 84 166 100
rect 170 92 174 100
rect 178 84 182 100
rect 186 84 190 92
rect 194 84 198 100
rect 204 94 208 98
rect 213 94 217 98
rect 222 94 226 98
rect 231 92 235 100
rect 239 92 243 100
rect 257 92 261 100
rect 274 92 278 100
rect 283 92 287 100
rect 293 92 297 100
<< m2contact >>
rect 45 113 50 118
rect 174 113 179 118
rect 9 59 14 64
rect 25 59 30 64
rect 69 65 74 70
rect 124 79 129 84
rect 117 56 122 61
rect 138 59 143 64
rect 154 59 159 64
rect 198 65 203 70
rect 53 10 58 15
rect 182 10 187 15
rect 269 5 274 10
<< psubstratepcontact >>
rect 2 20 6 24
rect 75 20 79 24
rect 93 20 97 24
rect 103 20 107 24
rect 131 20 135 24
rect 204 20 208 24
rect 222 20 226 24
rect 232 20 236 24
rect 265 20 269 24
rect 283 20 287 24
<< nsubstratencontact >>
rect 18 104 22 108
rect 76 104 80 108
rect 93 104 97 108
rect 147 104 151 108
rect 205 104 209 108
rect 222 104 226 108
rect 258 104 262 108
rect 283 104 287 108
<< labels >>
rlabel polycontact 4 82 4 82 3 A
rlabel polycontact 20 82 20 82 1 B
rlabel polycontact 149 82 149 82 1 C
rlabel metal1 299 85 299 85 7 carry
rlabel metal2 300 67 300 67 7 sum
rlabel metal1 119 106 119 106 1 VDD
rlabel metal1 115 22 115 22 1 GND
<< end >>
