* SPICE3 file created from /home/akhil/AND_GATE.ext - technology: scmos

.include bsim.txt
.option scale=0.09u
VDD vdd 0 DC 1.8
VA A 0 dc 1 pulse (0 1.8 190p 10p 10p 190p 400p)
VB B 0 dc 1 pulse (0 1.8 190p 10p 10p 190p 400p)

M1000 vout a_7_44# vdd Vdd pfet w=8 l=2
+  ad=40 pd=26 as=120 ps=78
M1001 a_7_44# A vdd Vdd pfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1002 vdd B a_7_44# Vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 vout a_7_44# Gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=60 ps=44
M1004 a_7_10# A Gnd Gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1005 a_7_44# B a_7_10# Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0

.tran 10p 2n
.control
run
set xbrushwidth = 2
plot A B+2 vout+4
.endc
.end

