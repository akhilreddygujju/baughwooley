magic
tech scmos
timestamp 1734110805
<< polysilicon >>
rect -1609 41 -1607 43
rect -1590 41 -1588 43
rect -1571 41 -1569 71
rect -1549 41 -1547 43
rect -1527 41 -1525 43
rect -1511 41 -1509 62
rect -1475 41 -1473 62
rect -1453 41 -1451 43
rect -1431 41 -1429 43
rect -1415 41 -1413 71
rect -1384 41 -1382 43
rect -1609 -2 -1607 33
rect -1590 -2 -1588 33
rect -1571 31 -1569 33
rect -1549 2 -1547 25
rect -1571 -2 -1569 0
rect -1527 -2 -1525 33
rect -1511 31 -1509 33
rect -1475 31 -1473 33
rect -1453 2 -1451 25
rect -1511 -2 -1509 0
rect -1475 -2 -1473 0
rect -1431 -2 -1429 33
rect -1415 31 -1413 33
rect -1415 -2 -1413 0
rect -1384 -2 -1382 33
rect -1609 -8 -1607 -6
rect -1590 -8 -1588 -6
rect -1571 -39 -1569 -6
rect -1549 -8 -1547 -6
rect -1527 -8 -1525 -6
rect -1511 -48 -1509 -6
rect -1475 -48 -1473 -6
rect -1453 -8 -1451 -6
rect -1431 -8 -1429 -6
rect -1415 -39 -1413 -6
rect -1384 -8 -1382 -6
rect -1611 -115 -1609 -113
rect -1592 -115 -1590 -113
rect -1573 -115 -1571 -85
rect -1551 -115 -1549 -113
rect -1529 -115 -1527 -113
rect -1513 -115 -1511 -94
rect -1477 -115 -1475 -94
rect -1455 -115 -1453 -113
rect -1433 -115 -1431 -113
rect -1417 -115 -1415 -85
rect -1386 -115 -1384 -113
rect -1611 -158 -1609 -123
rect -1592 -158 -1590 -123
rect -1573 -125 -1571 -123
rect -1551 -154 -1549 -131
rect -1573 -158 -1571 -156
rect -1529 -158 -1527 -123
rect -1513 -125 -1511 -123
rect -1477 -125 -1475 -123
rect -1455 -154 -1453 -131
rect -1513 -158 -1511 -156
rect -1477 -158 -1475 -156
rect -1433 -158 -1431 -123
rect -1417 -125 -1415 -123
rect -1417 -158 -1415 -156
rect -1386 -158 -1384 -123
rect -1611 -164 -1609 -162
rect -1592 -164 -1590 -162
rect -1573 -195 -1571 -162
rect -1551 -164 -1549 -162
rect -1529 -164 -1527 -162
rect -1513 -204 -1511 -162
rect -1477 -204 -1475 -162
rect -1455 -164 -1453 -162
rect -1433 -164 -1431 -162
rect -1417 -195 -1415 -162
rect -1386 -164 -1384 -162
rect -444 -205 -442 -179
rect -436 -205 -434 -179
rect -395 -192 -393 -179
rect -379 -192 -377 -138
rect -363 -192 -361 -179
rect -355 -192 -353 -190
rect -347 -192 -345 -179
rect -339 -192 -337 -190
rect -320 -192 -318 -180
rect -312 -192 -310 -180
rect -294 -192 -292 -190
rect -266 -192 -264 -179
rect -250 -192 -248 -138
rect -234 -192 -232 -179
rect -226 -192 -224 -190
rect -218 -192 -216 -179
rect -210 -192 -208 -190
rect -191 -192 -189 -180
rect -183 -192 -181 -180
rect -165 -192 -163 -190
rect -138 -192 -136 -180
rect -130 -192 -128 -180
rect -112 -192 -110 -190
rect -444 -239 -442 -213
rect -436 -239 -434 -213
rect -444 -249 -442 -247
rect -436 -249 -434 -247
rect -395 -260 -393 -200
rect -379 -260 -377 -200
rect -363 -256 -361 -208
rect -355 -256 -353 -208
rect -347 -256 -345 -208
rect -339 -256 -337 -208
rect -320 -256 -318 -200
rect -312 -256 -310 -200
rect -294 -260 -292 -200
rect -266 -260 -264 -200
rect -250 -260 -248 -200
rect -234 -256 -232 -208
rect -226 -256 -224 -208
rect -218 -256 -216 -208
rect -210 -256 -208 -208
rect -191 -256 -189 -200
rect -183 -256 -181 -200
rect -165 -260 -163 -200
rect -138 -255 -136 -200
rect -130 -255 -128 -200
rect -112 -260 -110 -200
rect -55 -208 -53 -179
rect -47 -208 -45 -179
rect 1 -192 3 -179
rect 17 -192 19 -161
rect 33 -192 35 -179
rect 41 -192 43 -190
rect 49 -192 51 -179
rect 57 -192 59 -190
rect 76 -192 78 -180
rect 84 -192 86 -180
rect 102 -192 104 -190
rect 130 -192 132 -179
rect 146 -192 148 -161
rect 162 -192 164 -179
rect 170 -192 172 -190
rect 178 -192 180 -179
rect 186 -192 188 -190
rect 205 -192 207 -180
rect 213 -192 215 -180
rect 231 -192 233 -190
rect 258 -192 260 -180
rect 266 -192 268 -180
rect 284 -192 286 -190
rect -31 -208 -29 -206
rect -55 -242 -53 -216
rect -47 -242 -45 -216
rect -31 -246 -29 -216
rect -55 -252 -53 -250
rect -47 -252 -45 -250
rect -31 -252 -29 -250
rect 1 -260 3 -200
rect 17 -260 19 -200
rect 33 -256 35 -208
rect 41 -256 43 -208
rect 49 -256 51 -208
rect 57 -256 59 -208
rect 76 -256 78 -200
rect 84 -256 86 -200
rect -395 -266 -393 -264
rect -379 -277 -377 -264
rect -363 -266 -361 -264
rect -355 -277 -353 -264
rect -347 -266 -345 -264
rect -339 -277 -337 -264
rect -320 -266 -318 -264
rect -312 -276 -310 -264
rect -294 -266 -292 -264
rect -266 -266 -264 -264
rect -250 -277 -248 -264
rect -234 -266 -232 -264
rect -226 -277 -224 -264
rect -218 -266 -216 -264
rect -210 -277 -208 -264
rect -191 -266 -189 -264
rect -183 -276 -181 -264
rect -165 -266 -163 -264
rect -138 -266 -136 -263
rect -130 -276 -128 -263
rect 102 -260 104 -200
rect 130 -260 132 -200
rect 146 -260 148 -200
rect 162 -256 164 -208
rect 170 -256 172 -208
rect 178 -256 180 -208
rect 186 -256 188 -208
rect 205 -256 207 -200
rect 213 -256 215 -200
rect 231 -260 233 -200
rect 258 -255 260 -200
rect 266 -255 268 -200
rect 284 -260 286 -200
rect -112 -266 -110 -264
rect 1 -266 3 -264
rect 17 -277 19 -264
rect 33 -266 35 -264
rect 41 -277 43 -264
rect 49 -266 51 -264
rect 57 -277 59 -264
rect 76 -266 78 -264
rect 84 -276 86 -264
rect 102 -266 104 -264
rect 130 -266 132 -264
rect 146 -277 148 -264
rect 162 -266 164 -264
rect 170 -277 172 -264
rect 178 -266 180 -264
rect 186 -277 188 -264
rect 205 -266 207 -264
rect 213 -276 215 -264
rect 231 -266 233 -264
rect 258 -266 260 -263
rect 266 -276 268 -263
rect 284 -266 286 -264
rect -1611 -323 -1609 -321
rect -1592 -323 -1590 -321
rect -1573 -323 -1571 -293
rect -1551 -323 -1549 -321
rect -1529 -323 -1527 -321
rect -1513 -323 -1511 -302
rect -1477 -323 -1475 -302
rect -1455 -323 -1453 -321
rect -1433 -323 -1431 -321
rect -1417 -323 -1415 -293
rect -1386 -323 -1384 -321
rect -1611 -366 -1609 -331
rect -1592 -366 -1590 -331
rect -1573 -333 -1571 -331
rect -1551 -362 -1549 -339
rect -1573 -366 -1571 -364
rect -1529 -366 -1527 -331
rect -1513 -333 -1511 -331
rect -1477 -333 -1475 -331
rect -1455 -362 -1453 -339
rect -1513 -366 -1511 -364
rect -1477 -366 -1475 -364
rect -1433 -366 -1431 -331
rect -1417 -333 -1415 -331
rect -1417 -366 -1415 -364
rect -1386 -366 -1384 -331
rect -422 -360 -420 -344
rect -659 -362 -420 -360
rect -385 -345 -250 -343
rect -1611 -372 -1609 -370
rect -1592 -372 -1590 -370
rect -1573 -403 -1571 -370
rect -1551 -372 -1549 -370
rect -1529 -372 -1527 -370
rect -1513 -412 -1511 -370
rect -1477 -412 -1475 -370
rect -1455 -372 -1453 -370
rect -1433 -372 -1431 -370
rect -1417 -403 -1415 -370
rect -1386 -372 -1384 -370
rect -860 -415 -858 -386
rect -852 -415 -850 -386
rect -804 -399 -802 -386
rect -788 -399 -786 -397
rect -772 -399 -770 -386
rect -764 -399 -762 -397
rect -756 -399 -754 -386
rect -748 -399 -746 -397
rect -729 -399 -727 -387
rect -721 -399 -719 -387
rect -703 -399 -701 -397
rect -675 -399 -673 -386
rect -659 -399 -657 -362
rect -643 -399 -641 -386
rect -635 -399 -633 -397
rect -627 -399 -625 -386
rect -619 -399 -617 -397
rect -600 -399 -598 -387
rect -592 -399 -590 -387
rect -574 -399 -572 -397
rect -547 -399 -545 -387
rect -539 -399 -537 -387
rect -521 -399 -519 -397
rect -836 -415 -834 -413
rect -860 -449 -858 -423
rect -852 -449 -850 -423
rect -836 -453 -834 -423
rect -860 -459 -858 -457
rect -852 -459 -850 -457
rect -836 -459 -834 -457
rect -804 -467 -802 -407
rect -788 -467 -786 -407
rect -772 -463 -770 -415
rect -764 -463 -762 -415
rect -756 -463 -754 -415
rect -748 -463 -746 -415
rect -729 -463 -727 -407
rect -721 -463 -719 -407
rect -703 -467 -701 -407
rect -675 -467 -673 -407
rect -659 -467 -657 -407
rect -643 -463 -641 -415
rect -635 -463 -633 -415
rect -627 -463 -625 -415
rect -619 -463 -617 -415
rect -600 -463 -598 -407
rect -592 -463 -590 -407
rect -574 -467 -572 -407
rect -547 -462 -545 -407
rect -539 -462 -537 -407
rect -521 -467 -519 -407
rect -450 -412 -448 -386
rect -442 -412 -440 -386
rect -401 -399 -399 -386
rect -385 -399 -383 -345
rect -256 -363 24 -361
rect -369 -399 -367 -386
rect -361 -399 -359 -397
rect -353 -399 -351 -386
rect -345 -399 -343 -397
rect -326 -399 -324 -387
rect -318 -399 -316 -387
rect -300 -399 -298 -397
rect -272 -399 -270 -386
rect -256 -399 -254 -363
rect -240 -399 -238 -386
rect -232 -399 -230 -397
rect -224 -399 -222 -386
rect -216 -399 -214 -397
rect -197 -399 -195 -387
rect -189 -399 -187 -387
rect -171 -399 -169 -397
rect -144 -399 -142 -387
rect -136 -399 -134 -387
rect -118 -399 -116 -397
rect -450 -446 -448 -420
rect -442 -446 -440 -420
rect -450 -456 -448 -454
rect -442 -456 -440 -454
rect -401 -467 -399 -407
rect -385 -467 -383 -407
rect -369 -463 -367 -415
rect -361 -463 -359 -415
rect -353 -463 -351 -415
rect -345 -463 -343 -415
rect -326 -463 -324 -407
rect -318 -463 -316 -407
rect -804 -473 -802 -471
rect -788 -484 -786 -471
rect -772 -473 -770 -471
rect -764 -484 -762 -471
rect -756 -473 -754 -471
rect -748 -484 -746 -471
rect -729 -473 -727 -471
rect -721 -483 -719 -471
rect -703 -473 -701 -471
rect -675 -473 -673 -471
rect -659 -484 -657 -471
rect -643 -473 -641 -471
rect -635 -484 -633 -471
rect -627 -473 -625 -471
rect -619 -484 -617 -471
rect -600 -473 -598 -471
rect -592 -483 -590 -471
rect -574 -473 -572 -471
rect -547 -473 -545 -470
rect -539 -483 -537 -470
rect -300 -467 -298 -407
rect -272 -467 -270 -407
rect -256 -467 -254 -407
rect -240 -463 -238 -415
rect -232 -463 -230 -415
rect -224 -463 -222 -415
rect -216 -463 -214 -415
rect -197 -463 -195 -407
rect -189 -463 -187 -407
rect -171 -467 -169 -407
rect -144 -462 -142 -407
rect -136 -462 -134 -407
rect -118 -467 -116 -407
rect -521 -473 -519 -471
rect -401 -473 -399 -471
rect -385 -484 -383 -471
rect -369 -473 -367 -471
rect -361 -484 -359 -471
rect -353 -473 -351 -471
rect -345 -484 -343 -471
rect -326 -473 -324 -471
rect -318 -483 -316 -471
rect -300 -473 -298 -471
rect -272 -473 -270 -471
rect -256 -484 -254 -471
rect -240 -473 -238 -471
rect -232 -484 -230 -471
rect -224 -473 -222 -471
rect -216 -484 -214 -471
rect -197 -473 -195 -471
rect -189 -483 -187 -471
rect -171 -473 -169 -471
rect -144 -473 -142 -470
rect -136 -483 -134 -470
rect -118 -473 -116 -471
rect -1614 -546 -1612 -544
rect -1595 -546 -1593 -544
rect -1576 -546 -1574 -516
rect -1554 -546 -1552 -544
rect -1532 -546 -1530 -544
rect -1516 -546 -1514 -525
rect -1480 -546 -1478 -525
rect -1458 -546 -1456 -544
rect -1436 -546 -1434 -544
rect -1420 -546 -1418 -516
rect -1389 -546 -1387 -544
rect -1614 -589 -1612 -554
rect -1595 -589 -1593 -554
rect -1576 -556 -1574 -554
rect -1554 -585 -1552 -562
rect -1576 -589 -1574 -587
rect -1532 -589 -1530 -554
rect -1516 -556 -1514 -554
rect -1480 -556 -1478 -554
rect -1458 -585 -1456 -562
rect -1516 -589 -1514 -587
rect -1480 -589 -1478 -587
rect -1436 -589 -1434 -554
rect -1420 -556 -1418 -554
rect -1420 -589 -1418 -587
rect -1389 -589 -1387 -554
rect -1614 -595 -1612 -593
rect -1595 -595 -1593 -593
rect -1576 -626 -1574 -593
rect -1554 -595 -1552 -593
rect -1532 -595 -1530 -593
rect -1516 -635 -1514 -593
rect -1480 -635 -1478 -593
rect -1458 -595 -1456 -593
rect -1436 -595 -1434 -593
rect -1420 -626 -1418 -593
rect -1389 -595 -1387 -593
rect -1229 -643 -1227 -630
rect -1213 -643 -1211 -566
rect -833 -603 -293 -601
rect -1197 -643 -1195 -630
rect -1189 -643 -1187 -641
rect -1181 -643 -1179 -630
rect -1173 -643 -1171 -641
rect -1154 -643 -1152 -631
rect -1146 -643 -1144 -631
rect -1128 -643 -1126 -641
rect -1100 -643 -1098 -630
rect -1084 -643 -1082 -604
rect -1068 -643 -1066 -630
rect -1060 -643 -1058 -641
rect -1052 -643 -1050 -630
rect -1044 -643 -1042 -641
rect -1025 -643 -1023 -631
rect -1017 -643 -1015 -631
rect -999 -643 -997 -641
rect -972 -643 -970 -631
rect -964 -643 -962 -631
rect -946 -643 -944 -641
rect -849 -643 -847 -630
rect -833 -643 -831 -603
rect -817 -643 -815 -630
rect -809 -643 -807 -641
rect -801 -643 -799 -630
rect -793 -643 -791 -641
rect -774 -643 -772 -631
rect -766 -643 -764 -631
rect -748 -643 -746 -641
rect -720 -643 -718 -630
rect -704 -643 -702 -641
rect -688 -643 -686 -630
rect -680 -643 -678 -641
rect -672 -643 -670 -630
rect -664 -643 -662 -641
rect -645 -643 -643 -631
rect -637 -643 -635 -631
rect -619 -643 -617 -641
rect -592 -643 -590 -631
rect -584 -643 -582 -631
rect -566 -643 -564 -641
rect -1229 -711 -1227 -651
rect -1213 -711 -1211 -651
rect -1197 -707 -1195 -659
rect -1189 -707 -1187 -659
rect -1181 -707 -1179 -659
rect -1173 -707 -1171 -659
rect -1154 -707 -1152 -651
rect -1146 -707 -1144 -651
rect -1128 -711 -1126 -651
rect -1100 -711 -1098 -651
rect -1084 -711 -1082 -651
rect -1068 -707 -1066 -659
rect -1060 -707 -1058 -659
rect -1052 -707 -1050 -659
rect -1044 -707 -1042 -659
rect -1025 -707 -1023 -651
rect -1017 -707 -1015 -651
rect -999 -711 -997 -651
rect -972 -706 -970 -651
rect -964 -706 -962 -651
rect -946 -711 -944 -651
rect -849 -711 -847 -651
rect -833 -711 -831 -651
rect -817 -707 -815 -659
rect -809 -707 -807 -659
rect -801 -707 -799 -659
rect -793 -707 -791 -659
rect -774 -707 -772 -651
rect -766 -707 -764 -651
rect -1229 -717 -1227 -715
rect -1213 -728 -1211 -715
rect -1197 -717 -1195 -715
rect -1189 -728 -1187 -715
rect -1181 -717 -1179 -715
rect -1173 -728 -1171 -715
rect -1154 -717 -1152 -715
rect -1146 -727 -1144 -715
rect -1128 -717 -1126 -715
rect -1100 -717 -1098 -715
rect -1084 -728 -1082 -715
rect -1068 -717 -1066 -715
rect -1060 -728 -1058 -715
rect -1052 -717 -1050 -715
rect -1044 -728 -1042 -715
rect -1025 -717 -1023 -715
rect -1017 -727 -1015 -715
rect -999 -717 -997 -715
rect -972 -717 -970 -714
rect -964 -727 -962 -714
rect -748 -711 -746 -651
rect -720 -711 -718 -651
rect -704 -711 -702 -651
rect -688 -707 -686 -659
rect -680 -707 -678 -659
rect -672 -707 -670 -659
rect -664 -707 -662 -659
rect -645 -707 -643 -651
rect -637 -707 -635 -651
rect -619 -711 -617 -651
rect -592 -706 -590 -651
rect -584 -706 -582 -651
rect -566 -711 -564 -651
rect -946 -717 -944 -715
rect -849 -717 -847 -715
rect -833 -728 -831 -715
rect -817 -717 -815 -715
rect -809 -728 -807 -715
rect -801 -717 -799 -715
rect -793 -728 -791 -715
rect -774 -717 -772 -715
rect -766 -727 -764 -715
rect -748 -717 -746 -715
rect -720 -717 -718 -715
rect -704 -728 -702 -715
rect -688 -717 -686 -715
rect -680 -728 -678 -715
rect -672 -717 -670 -715
rect -664 -728 -662 -715
rect -645 -717 -643 -715
rect -637 -727 -635 -715
rect -619 -717 -617 -715
rect -592 -717 -590 -714
rect -584 -727 -582 -714
rect -566 -717 -564 -715
rect -1195 -908 -1193 -906
rect -1176 -908 -1174 -816
rect -1157 -908 -1155 -878
rect -1135 -908 -1133 -906
rect -1113 -908 -1111 -906
rect -1097 -908 -1095 -887
rect -1061 -908 -1059 -887
rect -1039 -908 -1037 -906
rect -1017 -908 -1015 -906
rect -1001 -908 -999 -878
rect -805 -891 -803 -889
rect -786 -891 -784 -813
rect -294 -818 -276 -816
rect -767 -891 -765 -861
rect -745 -891 -743 -889
rect -723 -891 -721 -889
rect -707 -891 -705 -870
rect -671 -891 -669 -870
rect -649 -891 -647 -889
rect -627 -891 -625 -889
rect -611 -891 -609 -861
rect -580 -891 -578 -889
rect -313 -890 -311 -888
rect -294 -890 -292 -818
rect -275 -890 -273 -860
rect -253 -890 -251 -888
rect -231 -890 -229 -888
rect -215 -890 -213 -869
rect -179 -890 -177 -869
rect -157 -890 -155 -888
rect -135 -890 -133 -888
rect -119 -890 -117 -860
rect -88 -890 -86 -888
rect -970 -908 -968 -906
rect -1195 -951 -1193 -916
rect -1176 -951 -1174 -916
rect -1157 -918 -1155 -916
rect -1135 -947 -1133 -924
rect -1157 -951 -1155 -949
rect -1113 -951 -1111 -916
rect -1097 -918 -1095 -916
rect -1061 -918 -1059 -916
rect -1039 -947 -1037 -924
rect -1097 -951 -1095 -949
rect -1061 -951 -1059 -949
rect -1017 -951 -1015 -916
rect -1001 -918 -999 -916
rect -1001 -951 -999 -949
rect -970 -951 -968 -916
rect -805 -934 -803 -899
rect -786 -934 -784 -899
rect -767 -901 -765 -899
rect -745 -930 -743 -907
rect -767 -934 -765 -932
rect -723 -934 -721 -899
rect -707 -901 -705 -899
rect -671 -901 -669 -899
rect -649 -930 -647 -907
rect -707 -934 -705 -932
rect -671 -934 -669 -932
rect -627 -934 -625 -899
rect -611 -901 -609 -899
rect -611 -934 -609 -932
rect -580 -934 -578 -899
rect -313 -933 -311 -898
rect -294 -933 -292 -898
rect -275 -900 -273 -898
rect -253 -929 -251 -906
rect -275 -933 -273 -931
rect -231 -933 -229 -898
rect -215 -900 -213 -898
rect -179 -900 -177 -898
rect -157 -929 -155 -906
rect -215 -933 -213 -931
rect -179 -933 -177 -931
rect -135 -933 -133 -898
rect -119 -900 -117 -898
rect -119 -933 -117 -931
rect -88 -933 -86 -898
rect 98 -905 100 -903
rect 117 -905 119 -864
rect 136 -905 138 -875
rect 158 -905 160 -903
rect 180 -905 182 -903
rect 196 -905 198 -884
rect 232 -905 234 -884
rect 254 -905 256 -903
rect 276 -905 278 -903
rect 292 -905 294 -875
rect 323 -905 325 -903
rect -805 -940 -803 -938
rect -786 -940 -784 -938
rect -1195 -957 -1193 -955
rect -1176 -957 -1174 -955
rect -1157 -988 -1155 -955
rect -1135 -957 -1133 -955
rect -1113 -957 -1111 -955
rect -1097 -997 -1095 -955
rect -1061 -997 -1059 -955
rect -1039 -957 -1037 -955
rect -1017 -957 -1015 -955
rect -1001 -988 -999 -955
rect -970 -957 -968 -955
rect -767 -971 -765 -938
rect -745 -940 -743 -938
rect -723 -940 -721 -938
rect -707 -980 -705 -938
rect -671 -980 -669 -938
rect -649 -940 -647 -938
rect -627 -940 -625 -938
rect -611 -971 -609 -938
rect -580 -940 -578 -938
rect -313 -939 -311 -937
rect -294 -939 -292 -937
rect -275 -970 -273 -937
rect -253 -939 -251 -937
rect -231 -939 -229 -937
rect -215 -979 -213 -937
rect -179 -979 -177 -937
rect -157 -939 -155 -937
rect -135 -939 -133 -937
rect -119 -970 -117 -937
rect -88 -939 -86 -937
rect 98 -948 100 -913
rect 117 -948 119 -913
rect 136 -915 138 -913
rect 158 -944 160 -921
rect 136 -948 138 -946
rect 180 -948 182 -913
rect 196 -915 198 -913
rect 232 -915 234 -913
rect 254 -944 256 -921
rect 196 -948 198 -946
rect 232 -948 234 -946
rect 276 -948 278 -913
rect 292 -915 294 -913
rect 292 -948 294 -946
rect 323 -948 325 -913
rect 98 -954 100 -952
rect 117 -954 119 -952
rect 136 -985 138 -952
rect 158 -954 160 -952
rect 180 -954 182 -952
rect 196 -994 198 -952
rect 232 -994 234 -952
rect 254 -954 256 -952
rect 276 -954 278 -952
rect 292 -985 294 -952
rect 323 -954 325 -952
<< ndiffusion >>
rect -1610 -6 -1609 -2
rect -1607 -6 -1606 -2
rect -1591 -6 -1590 -2
rect -1588 -6 -1587 -2
rect -1572 -6 -1571 -2
rect -1569 -6 -1568 -2
rect -1550 -6 -1549 2
rect -1547 -6 -1546 2
rect -1528 -6 -1527 -2
rect -1525 -6 -1524 -2
rect -1512 -6 -1511 -2
rect -1509 -6 -1508 -2
rect -1476 -6 -1475 -2
rect -1473 -6 -1472 -2
rect -1454 -6 -1453 2
rect -1451 -6 -1450 2
rect -1432 -6 -1431 -2
rect -1429 -6 -1428 -2
rect -1416 -6 -1415 -2
rect -1413 -6 -1412 -2
rect -1385 -6 -1384 -2
rect -1382 -6 -1381 -2
rect -1612 -162 -1611 -158
rect -1609 -162 -1608 -158
rect -1593 -162 -1592 -158
rect -1590 -162 -1589 -158
rect -1574 -162 -1573 -158
rect -1571 -162 -1570 -158
rect -1552 -162 -1551 -154
rect -1549 -162 -1548 -154
rect -1530 -162 -1529 -158
rect -1527 -162 -1526 -158
rect -1514 -162 -1513 -158
rect -1511 -162 -1510 -158
rect -1478 -162 -1477 -158
rect -1475 -162 -1474 -158
rect -1456 -162 -1455 -154
rect -1453 -162 -1452 -154
rect -1434 -162 -1433 -158
rect -1431 -162 -1430 -158
rect -1418 -162 -1417 -158
rect -1415 -162 -1414 -158
rect -1387 -162 -1386 -158
rect -1384 -162 -1383 -158
rect -445 -247 -444 -239
rect -442 -247 -436 -239
rect -434 -247 -433 -239
rect -396 -264 -395 -260
rect -393 -264 -392 -260
rect -380 -264 -379 -260
rect -377 -264 -376 -260
rect -364 -264 -363 -256
rect -361 -264 -355 -256
rect -353 -264 -352 -256
rect -348 -264 -347 -256
rect -345 -264 -339 -256
rect -337 -264 -336 -256
rect -323 -264 -320 -256
rect -318 -264 -312 -256
rect -310 -264 -307 -256
rect -295 -264 -294 -260
rect -292 -264 -291 -260
rect -267 -264 -266 -260
rect -264 -264 -263 -260
rect -251 -264 -250 -260
rect -248 -264 -247 -260
rect -235 -264 -234 -256
rect -232 -264 -226 -256
rect -224 -264 -223 -256
rect -219 -264 -218 -256
rect -216 -264 -210 -256
rect -208 -264 -207 -256
rect -194 -264 -191 -256
rect -189 -264 -183 -256
rect -181 -264 -178 -256
rect -166 -264 -165 -260
rect -163 -264 -162 -260
rect -140 -263 -138 -255
rect -136 -263 -135 -255
rect -131 -263 -130 -255
rect -128 -263 -127 -255
rect -56 -250 -55 -242
rect -53 -250 -47 -242
rect -45 -250 -44 -242
rect -32 -250 -31 -246
rect -29 -250 -28 -246
rect -114 -264 -112 -260
rect -110 -264 -108 -260
rect 0 -264 1 -260
rect 3 -264 4 -260
rect 16 -264 17 -260
rect 19 -264 20 -260
rect 32 -264 33 -256
rect 35 -264 41 -256
rect 43 -264 44 -256
rect 48 -264 49 -256
rect 51 -264 57 -256
rect 59 -264 60 -256
rect 73 -264 76 -256
rect 78 -264 84 -256
rect 86 -264 89 -256
rect 101 -264 102 -260
rect 104 -264 105 -260
rect 129 -264 130 -260
rect 132 -264 133 -260
rect 145 -264 146 -260
rect 148 -264 149 -260
rect 161 -264 162 -256
rect 164 -264 170 -256
rect 172 -264 173 -256
rect 177 -264 178 -256
rect 180 -264 186 -256
rect 188 -264 189 -256
rect 202 -264 205 -256
rect 207 -264 213 -256
rect 215 -264 218 -256
rect 230 -264 231 -260
rect 233 -264 234 -260
rect 256 -263 258 -255
rect 260 -263 261 -255
rect 265 -263 266 -255
rect 268 -263 269 -255
rect 282 -264 284 -260
rect 286 -264 288 -260
rect -1612 -370 -1611 -366
rect -1609 -370 -1608 -366
rect -1593 -370 -1592 -366
rect -1590 -370 -1589 -366
rect -1574 -370 -1573 -366
rect -1571 -370 -1570 -366
rect -1552 -370 -1551 -362
rect -1549 -370 -1548 -362
rect -1530 -370 -1529 -366
rect -1527 -370 -1526 -366
rect -1514 -370 -1513 -366
rect -1511 -370 -1510 -366
rect -1478 -370 -1477 -366
rect -1475 -370 -1474 -366
rect -1456 -370 -1455 -362
rect -1453 -370 -1452 -362
rect -1434 -370 -1433 -366
rect -1431 -370 -1430 -366
rect -1418 -370 -1417 -366
rect -1415 -370 -1414 -366
rect -1387 -370 -1386 -366
rect -1384 -370 -1383 -366
rect -861 -457 -860 -449
rect -858 -457 -852 -449
rect -850 -457 -849 -449
rect -837 -457 -836 -453
rect -834 -457 -833 -453
rect -805 -471 -804 -467
rect -802 -471 -801 -467
rect -789 -471 -788 -467
rect -786 -471 -785 -467
rect -773 -471 -772 -463
rect -770 -471 -764 -463
rect -762 -471 -761 -463
rect -757 -471 -756 -463
rect -754 -471 -748 -463
rect -746 -471 -745 -463
rect -732 -471 -729 -463
rect -727 -471 -721 -463
rect -719 -471 -716 -463
rect -704 -471 -703 -467
rect -701 -471 -700 -467
rect -676 -471 -675 -467
rect -673 -471 -672 -467
rect -660 -471 -659 -467
rect -657 -471 -656 -467
rect -644 -471 -643 -463
rect -641 -471 -635 -463
rect -633 -471 -632 -463
rect -628 -471 -627 -463
rect -625 -471 -619 -463
rect -617 -471 -616 -463
rect -603 -471 -600 -463
rect -598 -471 -592 -463
rect -590 -471 -587 -463
rect -575 -471 -574 -467
rect -572 -471 -571 -467
rect -549 -470 -547 -462
rect -545 -470 -544 -462
rect -540 -470 -539 -462
rect -537 -470 -536 -462
rect -451 -454 -450 -446
rect -448 -454 -442 -446
rect -440 -454 -439 -446
rect -523 -471 -521 -467
rect -519 -471 -517 -467
rect -402 -471 -401 -467
rect -399 -471 -398 -467
rect -386 -471 -385 -467
rect -383 -471 -382 -467
rect -370 -471 -369 -463
rect -367 -471 -361 -463
rect -359 -471 -358 -463
rect -354 -471 -353 -463
rect -351 -471 -345 -463
rect -343 -471 -342 -463
rect -329 -471 -326 -463
rect -324 -471 -318 -463
rect -316 -471 -313 -463
rect -301 -471 -300 -467
rect -298 -471 -297 -467
rect -273 -471 -272 -467
rect -270 -471 -269 -467
rect -257 -471 -256 -467
rect -254 -471 -253 -467
rect -241 -471 -240 -463
rect -238 -471 -232 -463
rect -230 -471 -229 -463
rect -225 -471 -224 -463
rect -222 -471 -216 -463
rect -214 -471 -213 -463
rect -200 -471 -197 -463
rect -195 -471 -189 -463
rect -187 -471 -184 -463
rect -172 -471 -171 -467
rect -169 -471 -168 -467
rect -146 -470 -144 -462
rect -142 -470 -141 -462
rect -137 -470 -136 -462
rect -134 -470 -133 -462
rect -120 -471 -118 -467
rect -116 -471 -114 -467
rect -1615 -593 -1614 -589
rect -1612 -593 -1611 -589
rect -1596 -593 -1595 -589
rect -1593 -593 -1592 -589
rect -1577 -593 -1576 -589
rect -1574 -593 -1573 -589
rect -1555 -593 -1554 -585
rect -1552 -593 -1551 -585
rect -1533 -593 -1532 -589
rect -1530 -593 -1529 -589
rect -1517 -593 -1516 -589
rect -1514 -593 -1513 -589
rect -1481 -593 -1480 -589
rect -1478 -593 -1477 -589
rect -1459 -593 -1458 -585
rect -1456 -593 -1455 -585
rect -1437 -593 -1436 -589
rect -1434 -593 -1433 -589
rect -1421 -593 -1420 -589
rect -1418 -593 -1417 -589
rect -1390 -593 -1389 -589
rect -1387 -593 -1386 -589
rect -1230 -715 -1229 -711
rect -1227 -715 -1226 -711
rect -1214 -715 -1213 -711
rect -1211 -715 -1210 -711
rect -1198 -715 -1197 -707
rect -1195 -715 -1189 -707
rect -1187 -715 -1186 -707
rect -1182 -715 -1181 -707
rect -1179 -715 -1173 -707
rect -1171 -715 -1170 -707
rect -1157 -715 -1154 -707
rect -1152 -715 -1146 -707
rect -1144 -715 -1141 -707
rect -1129 -715 -1128 -711
rect -1126 -715 -1125 -711
rect -1101 -715 -1100 -711
rect -1098 -715 -1097 -711
rect -1085 -715 -1084 -711
rect -1082 -715 -1081 -711
rect -1069 -715 -1068 -707
rect -1066 -715 -1060 -707
rect -1058 -715 -1057 -707
rect -1053 -715 -1052 -707
rect -1050 -715 -1044 -707
rect -1042 -715 -1041 -707
rect -1028 -715 -1025 -707
rect -1023 -715 -1017 -707
rect -1015 -715 -1012 -707
rect -1000 -715 -999 -711
rect -997 -715 -996 -711
rect -974 -714 -972 -706
rect -970 -714 -969 -706
rect -965 -714 -964 -706
rect -962 -714 -961 -706
rect -948 -715 -946 -711
rect -944 -715 -942 -711
rect -850 -715 -849 -711
rect -847 -715 -846 -711
rect -834 -715 -833 -711
rect -831 -715 -830 -711
rect -818 -715 -817 -707
rect -815 -715 -809 -707
rect -807 -715 -806 -707
rect -802 -715 -801 -707
rect -799 -715 -793 -707
rect -791 -715 -790 -707
rect -777 -715 -774 -707
rect -772 -715 -766 -707
rect -764 -715 -761 -707
rect -749 -715 -748 -711
rect -746 -715 -745 -711
rect -721 -715 -720 -711
rect -718 -715 -717 -711
rect -705 -715 -704 -711
rect -702 -715 -701 -711
rect -689 -715 -688 -707
rect -686 -715 -680 -707
rect -678 -715 -677 -707
rect -673 -715 -672 -707
rect -670 -715 -664 -707
rect -662 -715 -661 -707
rect -648 -715 -645 -707
rect -643 -715 -637 -707
rect -635 -715 -632 -707
rect -620 -715 -619 -711
rect -617 -715 -616 -711
rect -594 -714 -592 -706
rect -590 -714 -589 -706
rect -585 -714 -584 -706
rect -582 -714 -581 -706
rect -568 -715 -566 -711
rect -564 -715 -562 -711
rect -1196 -955 -1195 -951
rect -1193 -955 -1192 -951
rect -1177 -955 -1176 -951
rect -1174 -955 -1173 -951
rect -1158 -955 -1157 -951
rect -1155 -955 -1154 -951
rect -1136 -955 -1135 -947
rect -1133 -955 -1132 -947
rect -1114 -955 -1113 -951
rect -1111 -955 -1110 -951
rect -1098 -955 -1097 -951
rect -1095 -955 -1094 -951
rect -1062 -955 -1061 -951
rect -1059 -955 -1058 -951
rect -1040 -955 -1039 -947
rect -1037 -955 -1036 -947
rect -806 -938 -805 -934
rect -803 -938 -802 -934
rect -787 -938 -786 -934
rect -784 -938 -783 -934
rect -768 -938 -767 -934
rect -765 -938 -764 -934
rect -746 -938 -745 -930
rect -743 -938 -742 -930
rect -724 -938 -723 -934
rect -721 -938 -720 -934
rect -708 -938 -707 -934
rect -705 -938 -704 -934
rect -672 -938 -671 -934
rect -669 -938 -668 -934
rect -650 -938 -649 -930
rect -647 -938 -646 -930
rect -628 -938 -627 -934
rect -625 -938 -624 -934
rect -612 -938 -611 -934
rect -609 -938 -608 -934
rect -581 -938 -580 -934
rect -578 -938 -577 -934
rect -314 -937 -313 -933
rect -311 -937 -310 -933
rect -295 -937 -294 -933
rect -292 -937 -291 -933
rect -276 -937 -275 -933
rect -273 -937 -272 -933
rect -254 -937 -253 -929
rect -251 -937 -250 -929
rect -232 -937 -231 -933
rect -229 -937 -228 -933
rect -216 -937 -215 -933
rect -213 -937 -212 -933
rect -180 -937 -179 -933
rect -177 -937 -176 -933
rect -158 -937 -157 -929
rect -155 -937 -154 -929
rect -136 -937 -135 -933
rect -133 -937 -132 -933
rect -120 -937 -119 -933
rect -117 -937 -116 -933
rect -89 -937 -88 -933
rect -86 -937 -85 -933
rect -1018 -955 -1017 -951
rect -1015 -955 -1014 -951
rect -1002 -955 -1001 -951
rect -999 -955 -998 -951
rect -971 -955 -970 -951
rect -968 -955 -967 -951
rect 97 -952 98 -948
rect 100 -952 101 -948
rect 116 -952 117 -948
rect 119 -952 120 -948
rect 135 -952 136 -948
rect 138 -952 139 -948
rect 157 -952 158 -944
rect 160 -952 161 -944
rect 179 -952 180 -948
rect 182 -952 183 -948
rect 195 -952 196 -948
rect 198 -952 199 -948
rect 231 -952 232 -948
rect 234 -952 235 -948
rect 253 -952 254 -944
rect 256 -952 257 -944
rect 275 -952 276 -948
rect 278 -952 279 -948
rect 291 -952 292 -948
rect 294 -952 295 -948
rect 322 -952 323 -948
rect 325 -952 326 -948
<< pdiffusion >>
rect -1610 33 -1609 41
rect -1607 33 -1606 41
rect -1591 33 -1590 41
rect -1588 33 -1587 41
rect -1572 33 -1571 41
rect -1569 33 -1568 41
rect -1550 25 -1549 41
rect -1547 25 -1546 41
rect -1528 33 -1527 41
rect -1525 33 -1524 41
rect -1512 33 -1511 41
rect -1509 33 -1508 41
rect -1476 33 -1475 41
rect -1473 33 -1472 41
rect -1454 25 -1453 41
rect -1451 25 -1450 41
rect -1432 33 -1431 41
rect -1429 33 -1428 41
rect -1416 33 -1415 41
rect -1413 33 -1412 41
rect -1385 33 -1384 41
rect -1382 33 -1381 41
rect -1612 -123 -1611 -115
rect -1609 -123 -1608 -115
rect -1593 -123 -1592 -115
rect -1590 -123 -1589 -115
rect -1574 -123 -1573 -115
rect -1571 -123 -1570 -115
rect -1552 -131 -1551 -115
rect -1549 -131 -1548 -115
rect -1530 -123 -1529 -115
rect -1527 -123 -1526 -115
rect -1514 -123 -1513 -115
rect -1511 -123 -1510 -115
rect -1478 -123 -1477 -115
rect -1475 -123 -1474 -115
rect -1456 -131 -1455 -115
rect -1453 -131 -1452 -115
rect -1434 -123 -1433 -115
rect -1431 -123 -1430 -115
rect -1418 -123 -1417 -115
rect -1415 -123 -1414 -115
rect -1387 -123 -1386 -115
rect -1384 -123 -1383 -115
rect -396 -200 -395 -192
rect -393 -200 -392 -192
rect -380 -200 -379 -192
rect -377 -200 -376 -192
rect -445 -213 -444 -205
rect -442 -213 -441 -205
rect -437 -213 -436 -205
rect -434 -213 -433 -205
rect -364 -208 -363 -192
rect -361 -200 -360 -192
rect -356 -200 -355 -192
rect -361 -208 -355 -200
rect -353 -208 -352 -192
rect -348 -208 -347 -192
rect -345 -200 -339 -192
rect -345 -208 -344 -200
rect -340 -208 -339 -200
rect -337 -208 -336 -192
rect -327 -194 -320 -192
rect -327 -198 -326 -194
rect -322 -198 -320 -194
rect -327 -200 -320 -198
rect -318 -194 -312 -192
rect -318 -198 -317 -194
rect -313 -198 -312 -194
rect -318 -200 -312 -198
rect -310 -194 -303 -192
rect -310 -198 -308 -194
rect -304 -198 -303 -194
rect -310 -200 -303 -198
rect -295 -200 -294 -192
rect -292 -200 -291 -192
rect -267 -200 -266 -192
rect -264 -200 -263 -192
rect -251 -200 -250 -192
rect -248 -200 -247 -192
rect -235 -208 -234 -192
rect -232 -200 -231 -192
rect -227 -200 -226 -192
rect -232 -208 -226 -200
rect -224 -208 -223 -192
rect -219 -208 -218 -192
rect -216 -200 -210 -192
rect -216 -208 -215 -200
rect -211 -208 -210 -200
rect -208 -208 -207 -192
rect -198 -194 -191 -192
rect -198 -198 -197 -194
rect -193 -198 -191 -194
rect -198 -200 -191 -198
rect -189 -194 -183 -192
rect -189 -198 -188 -194
rect -184 -198 -183 -194
rect -189 -200 -183 -198
rect -181 -194 -174 -192
rect -181 -198 -179 -194
rect -175 -198 -174 -194
rect -181 -200 -174 -198
rect -166 -200 -165 -192
rect -163 -200 -162 -192
rect -140 -200 -138 -192
rect -136 -200 -130 -192
rect -128 -200 -127 -192
rect -114 -200 -112 -192
rect -110 -200 -108 -192
rect 0 -200 1 -192
rect 3 -200 4 -192
rect 16 -200 17 -192
rect 19 -200 20 -192
rect -56 -216 -55 -208
rect -53 -216 -52 -208
rect -48 -216 -47 -208
rect -45 -216 -44 -208
rect -32 -216 -31 -208
rect -29 -216 -28 -208
rect 32 -208 33 -192
rect 35 -200 36 -192
rect 40 -200 41 -192
rect 35 -208 41 -200
rect 43 -208 44 -192
rect 48 -208 49 -192
rect 51 -200 57 -192
rect 51 -208 52 -200
rect 56 -208 57 -200
rect 59 -208 60 -192
rect 69 -194 76 -192
rect 69 -198 70 -194
rect 74 -198 76 -194
rect 69 -200 76 -198
rect 78 -194 84 -192
rect 78 -198 79 -194
rect 83 -198 84 -194
rect 78 -200 84 -198
rect 86 -194 93 -192
rect 86 -198 88 -194
rect 92 -198 93 -194
rect 86 -200 93 -198
rect 101 -200 102 -192
rect 104 -200 105 -192
rect 129 -200 130 -192
rect 132 -200 133 -192
rect 145 -200 146 -192
rect 148 -200 149 -192
rect 161 -208 162 -192
rect 164 -200 165 -192
rect 169 -200 170 -192
rect 164 -208 170 -200
rect 172 -208 173 -192
rect 177 -208 178 -192
rect 180 -200 186 -192
rect 180 -208 181 -200
rect 185 -208 186 -200
rect 188 -208 189 -192
rect 198 -194 205 -192
rect 198 -198 199 -194
rect 203 -198 205 -194
rect 198 -200 205 -198
rect 207 -194 213 -192
rect 207 -198 208 -194
rect 212 -198 213 -194
rect 207 -200 213 -198
rect 215 -194 222 -192
rect 215 -198 217 -194
rect 221 -198 222 -194
rect 215 -200 222 -198
rect 230 -200 231 -192
rect 233 -200 234 -192
rect 256 -200 258 -192
rect 260 -200 266 -192
rect 268 -200 269 -192
rect 282 -200 284 -192
rect 286 -200 288 -192
rect -1612 -331 -1611 -323
rect -1609 -331 -1608 -323
rect -1593 -331 -1592 -323
rect -1590 -331 -1589 -323
rect -1574 -331 -1573 -323
rect -1571 -331 -1570 -323
rect -1552 -339 -1551 -323
rect -1549 -339 -1548 -323
rect -1530 -331 -1529 -323
rect -1527 -331 -1526 -323
rect -1514 -331 -1513 -323
rect -1511 -331 -1510 -323
rect -1478 -331 -1477 -323
rect -1475 -331 -1474 -323
rect -1456 -339 -1455 -323
rect -1453 -339 -1452 -323
rect -1434 -331 -1433 -323
rect -1431 -331 -1430 -323
rect -1418 -331 -1417 -323
rect -1415 -331 -1414 -323
rect -1387 -331 -1386 -323
rect -1384 -331 -1383 -323
rect -805 -407 -804 -399
rect -802 -407 -801 -399
rect -789 -407 -788 -399
rect -786 -407 -785 -399
rect -861 -423 -860 -415
rect -858 -423 -857 -415
rect -853 -423 -852 -415
rect -850 -423 -849 -415
rect -837 -423 -836 -415
rect -834 -423 -833 -415
rect -773 -415 -772 -399
rect -770 -407 -769 -399
rect -765 -407 -764 -399
rect -770 -415 -764 -407
rect -762 -415 -761 -399
rect -757 -415 -756 -399
rect -754 -407 -748 -399
rect -754 -415 -753 -407
rect -749 -415 -748 -407
rect -746 -415 -745 -399
rect -736 -401 -729 -399
rect -736 -405 -735 -401
rect -731 -405 -729 -401
rect -736 -407 -729 -405
rect -727 -401 -721 -399
rect -727 -405 -726 -401
rect -722 -405 -721 -401
rect -727 -407 -721 -405
rect -719 -401 -712 -399
rect -719 -405 -717 -401
rect -713 -405 -712 -401
rect -719 -407 -712 -405
rect -704 -407 -703 -399
rect -701 -407 -700 -399
rect -676 -407 -675 -399
rect -673 -407 -672 -399
rect -660 -407 -659 -399
rect -657 -407 -656 -399
rect -644 -415 -643 -399
rect -641 -407 -640 -399
rect -636 -407 -635 -399
rect -641 -415 -635 -407
rect -633 -415 -632 -399
rect -628 -415 -627 -399
rect -625 -407 -619 -399
rect -625 -415 -624 -407
rect -620 -415 -619 -407
rect -617 -415 -616 -399
rect -607 -401 -600 -399
rect -607 -405 -606 -401
rect -602 -405 -600 -401
rect -607 -407 -600 -405
rect -598 -401 -592 -399
rect -598 -405 -597 -401
rect -593 -405 -592 -401
rect -598 -407 -592 -405
rect -590 -401 -583 -399
rect -590 -405 -588 -401
rect -584 -405 -583 -401
rect -590 -407 -583 -405
rect -575 -407 -574 -399
rect -572 -407 -571 -399
rect -549 -407 -547 -399
rect -545 -407 -539 -399
rect -537 -407 -536 -399
rect -523 -407 -521 -399
rect -519 -407 -517 -399
rect -402 -407 -401 -399
rect -399 -407 -398 -399
rect -386 -407 -385 -399
rect -383 -407 -382 -399
rect -451 -420 -450 -412
rect -448 -420 -447 -412
rect -443 -420 -442 -412
rect -440 -420 -439 -412
rect -370 -415 -369 -399
rect -367 -407 -366 -399
rect -362 -407 -361 -399
rect -367 -415 -361 -407
rect -359 -415 -358 -399
rect -354 -415 -353 -399
rect -351 -407 -345 -399
rect -351 -415 -350 -407
rect -346 -415 -345 -407
rect -343 -415 -342 -399
rect -333 -401 -326 -399
rect -333 -405 -332 -401
rect -328 -405 -326 -401
rect -333 -407 -326 -405
rect -324 -401 -318 -399
rect -324 -405 -323 -401
rect -319 -405 -318 -401
rect -324 -407 -318 -405
rect -316 -401 -309 -399
rect -316 -405 -314 -401
rect -310 -405 -309 -401
rect -316 -407 -309 -405
rect -301 -407 -300 -399
rect -298 -407 -297 -399
rect -273 -407 -272 -399
rect -270 -407 -269 -399
rect -257 -407 -256 -399
rect -254 -407 -253 -399
rect -241 -415 -240 -399
rect -238 -407 -237 -399
rect -233 -407 -232 -399
rect -238 -415 -232 -407
rect -230 -415 -229 -399
rect -225 -415 -224 -399
rect -222 -407 -216 -399
rect -222 -415 -221 -407
rect -217 -415 -216 -407
rect -214 -415 -213 -399
rect -204 -401 -197 -399
rect -204 -405 -203 -401
rect -199 -405 -197 -401
rect -204 -407 -197 -405
rect -195 -401 -189 -399
rect -195 -405 -194 -401
rect -190 -405 -189 -401
rect -195 -407 -189 -405
rect -187 -401 -180 -399
rect -187 -405 -185 -401
rect -181 -405 -180 -401
rect -187 -407 -180 -405
rect -172 -407 -171 -399
rect -169 -407 -168 -399
rect -146 -407 -144 -399
rect -142 -407 -136 -399
rect -134 -407 -133 -399
rect -120 -407 -118 -399
rect -116 -407 -114 -399
rect -1615 -554 -1614 -546
rect -1612 -554 -1611 -546
rect -1596 -554 -1595 -546
rect -1593 -554 -1592 -546
rect -1577 -554 -1576 -546
rect -1574 -554 -1573 -546
rect -1555 -562 -1554 -546
rect -1552 -562 -1551 -546
rect -1533 -554 -1532 -546
rect -1530 -554 -1529 -546
rect -1517 -554 -1516 -546
rect -1514 -554 -1513 -546
rect -1481 -554 -1480 -546
rect -1478 -554 -1477 -546
rect -1459 -562 -1458 -546
rect -1456 -562 -1455 -546
rect -1437 -554 -1436 -546
rect -1434 -554 -1433 -546
rect -1421 -554 -1420 -546
rect -1418 -554 -1417 -546
rect -1390 -554 -1389 -546
rect -1387 -554 -1386 -546
rect -1230 -651 -1229 -643
rect -1227 -651 -1226 -643
rect -1214 -651 -1213 -643
rect -1211 -651 -1210 -643
rect -1198 -659 -1197 -643
rect -1195 -651 -1194 -643
rect -1190 -651 -1189 -643
rect -1195 -659 -1189 -651
rect -1187 -659 -1186 -643
rect -1182 -659 -1181 -643
rect -1179 -651 -1173 -643
rect -1179 -659 -1178 -651
rect -1174 -659 -1173 -651
rect -1171 -659 -1170 -643
rect -1161 -645 -1154 -643
rect -1161 -649 -1160 -645
rect -1156 -649 -1154 -645
rect -1161 -651 -1154 -649
rect -1152 -645 -1146 -643
rect -1152 -649 -1151 -645
rect -1147 -649 -1146 -645
rect -1152 -651 -1146 -649
rect -1144 -645 -1137 -643
rect -1144 -649 -1142 -645
rect -1138 -649 -1137 -645
rect -1144 -651 -1137 -649
rect -1129 -651 -1128 -643
rect -1126 -651 -1125 -643
rect -1101 -651 -1100 -643
rect -1098 -651 -1097 -643
rect -1085 -651 -1084 -643
rect -1082 -651 -1081 -643
rect -1069 -659 -1068 -643
rect -1066 -651 -1065 -643
rect -1061 -651 -1060 -643
rect -1066 -659 -1060 -651
rect -1058 -659 -1057 -643
rect -1053 -659 -1052 -643
rect -1050 -651 -1044 -643
rect -1050 -659 -1049 -651
rect -1045 -659 -1044 -651
rect -1042 -659 -1041 -643
rect -1032 -645 -1025 -643
rect -1032 -649 -1031 -645
rect -1027 -649 -1025 -645
rect -1032 -651 -1025 -649
rect -1023 -645 -1017 -643
rect -1023 -649 -1022 -645
rect -1018 -649 -1017 -645
rect -1023 -651 -1017 -649
rect -1015 -645 -1008 -643
rect -1015 -649 -1013 -645
rect -1009 -649 -1008 -645
rect -1015 -651 -1008 -649
rect -1000 -651 -999 -643
rect -997 -651 -996 -643
rect -974 -651 -972 -643
rect -970 -651 -964 -643
rect -962 -651 -961 -643
rect -948 -651 -946 -643
rect -944 -651 -942 -643
rect -850 -651 -849 -643
rect -847 -651 -846 -643
rect -834 -651 -833 -643
rect -831 -651 -830 -643
rect -818 -659 -817 -643
rect -815 -651 -814 -643
rect -810 -651 -809 -643
rect -815 -659 -809 -651
rect -807 -659 -806 -643
rect -802 -659 -801 -643
rect -799 -651 -793 -643
rect -799 -659 -798 -651
rect -794 -659 -793 -651
rect -791 -659 -790 -643
rect -781 -645 -774 -643
rect -781 -649 -780 -645
rect -776 -649 -774 -645
rect -781 -651 -774 -649
rect -772 -645 -766 -643
rect -772 -649 -771 -645
rect -767 -649 -766 -645
rect -772 -651 -766 -649
rect -764 -645 -757 -643
rect -764 -649 -762 -645
rect -758 -649 -757 -645
rect -764 -651 -757 -649
rect -749 -651 -748 -643
rect -746 -651 -745 -643
rect -721 -651 -720 -643
rect -718 -651 -717 -643
rect -705 -651 -704 -643
rect -702 -651 -701 -643
rect -689 -659 -688 -643
rect -686 -651 -685 -643
rect -681 -651 -680 -643
rect -686 -659 -680 -651
rect -678 -659 -677 -643
rect -673 -659 -672 -643
rect -670 -651 -664 -643
rect -670 -659 -669 -651
rect -665 -659 -664 -651
rect -662 -659 -661 -643
rect -652 -645 -645 -643
rect -652 -649 -651 -645
rect -647 -649 -645 -645
rect -652 -651 -645 -649
rect -643 -645 -637 -643
rect -643 -649 -642 -645
rect -638 -649 -637 -645
rect -643 -651 -637 -649
rect -635 -645 -628 -643
rect -635 -649 -633 -645
rect -629 -649 -628 -645
rect -635 -651 -628 -649
rect -620 -651 -619 -643
rect -617 -651 -616 -643
rect -594 -651 -592 -643
rect -590 -651 -584 -643
rect -582 -651 -581 -643
rect -568 -651 -566 -643
rect -564 -651 -562 -643
rect -806 -899 -805 -891
rect -803 -899 -802 -891
rect -787 -899 -786 -891
rect -784 -899 -783 -891
rect -768 -899 -767 -891
rect -765 -899 -764 -891
rect -1196 -916 -1195 -908
rect -1193 -916 -1192 -908
rect -1177 -916 -1176 -908
rect -1174 -916 -1173 -908
rect -1158 -916 -1157 -908
rect -1155 -916 -1154 -908
rect -1136 -924 -1135 -908
rect -1133 -924 -1132 -908
rect -1114 -916 -1113 -908
rect -1111 -916 -1110 -908
rect -1098 -916 -1097 -908
rect -1095 -916 -1094 -908
rect -1062 -916 -1061 -908
rect -1059 -916 -1058 -908
rect -1040 -924 -1039 -908
rect -1037 -924 -1036 -908
rect -1018 -916 -1017 -908
rect -1015 -916 -1014 -908
rect -1002 -916 -1001 -908
rect -999 -916 -998 -908
rect -971 -916 -970 -908
rect -968 -916 -967 -908
rect -746 -907 -745 -891
rect -743 -907 -742 -891
rect -724 -899 -723 -891
rect -721 -899 -720 -891
rect -708 -899 -707 -891
rect -705 -899 -704 -891
rect -672 -899 -671 -891
rect -669 -899 -668 -891
rect -650 -907 -649 -891
rect -647 -907 -646 -891
rect -628 -899 -627 -891
rect -625 -899 -624 -891
rect -612 -899 -611 -891
rect -609 -899 -608 -891
rect -581 -899 -580 -891
rect -578 -899 -577 -891
rect -314 -898 -313 -890
rect -311 -898 -310 -890
rect -295 -898 -294 -890
rect -292 -898 -291 -890
rect -276 -898 -275 -890
rect -273 -898 -272 -890
rect -254 -906 -253 -890
rect -251 -906 -250 -890
rect -232 -898 -231 -890
rect -229 -898 -228 -890
rect -216 -898 -215 -890
rect -213 -898 -212 -890
rect -180 -898 -179 -890
rect -177 -898 -176 -890
rect -158 -906 -157 -890
rect -155 -906 -154 -890
rect -136 -898 -135 -890
rect -133 -898 -132 -890
rect -120 -898 -119 -890
rect -117 -898 -116 -890
rect -89 -898 -88 -890
rect -86 -898 -85 -890
rect 97 -913 98 -905
rect 100 -913 101 -905
rect 116 -913 117 -905
rect 119 -913 120 -905
rect 135 -913 136 -905
rect 138 -913 139 -905
rect 157 -921 158 -905
rect 160 -921 161 -905
rect 179 -913 180 -905
rect 182 -913 183 -905
rect 195 -913 196 -905
rect 198 -913 199 -905
rect 231 -913 232 -905
rect 234 -913 235 -905
rect 253 -921 254 -905
rect 256 -921 257 -905
rect 275 -913 276 -905
rect 278 -913 279 -905
rect 291 -913 292 -905
rect 294 -913 295 -905
rect 322 -913 323 -905
rect 325 -913 326 -905
<< metal1 >>
rect -1733 -64 -1724 127
rect -1625 106 378 123
rect -1624 71 -1572 75
rect -1568 71 -1416 75
rect -1624 17 -1620 71
rect -1600 62 -1512 66
rect -1508 62 -1476 66
rect -1354 50 -1349 106
rect -1614 49 -1349 50
rect -1614 45 -1613 49
rect -1609 45 -1594 49
rect -1590 45 -1553 49
rect -1549 45 -1531 49
rect -1527 45 -1457 49
rect -1453 45 -1435 49
rect -1431 45 -1388 49
rect -1384 45 -1349 49
rect -1614 44 -1349 45
rect -1614 41 -1610 44
rect -1595 41 -1591 44
rect -1554 41 -1550 44
rect -1532 41 -1528 44
rect -1458 41 -1454 44
rect -1436 41 -1432 44
rect -1389 41 -1385 44
rect -1606 18 -1602 33
rect -1624 13 -1613 17
rect -1587 17 -1583 33
rect -1576 17 -1572 33
rect -1587 13 -1572 17
rect -1624 -48 -1620 13
rect -1606 -2 -1602 13
rect -1587 -2 -1583 13
rect -1576 -2 -1572 13
rect -1568 18 -1564 33
rect -1546 17 -1542 25
rect -1524 17 -1520 33
rect -1516 17 -1512 33
rect -1563 13 -1553 17
rect -1546 13 -1539 17
rect -1535 13 -1531 17
rect -1524 13 -1512 17
rect -1568 -2 -1564 13
rect -1546 2 -1542 13
rect -1524 -2 -1520 13
rect -1516 -2 -1512 13
rect -1508 18 -1504 33
rect -1480 18 -1476 33
rect -1508 -2 -1504 13
rect -1480 -2 -1476 13
rect -1472 17 -1468 33
rect -1472 13 -1464 17
rect -1450 17 -1446 25
rect -1459 13 -1457 17
rect -1450 13 -1443 17
rect -1428 17 -1424 33
rect -1420 17 -1416 33
rect -1438 13 -1435 17
rect -1428 13 -1416 17
rect -1472 -2 -1468 13
rect -1450 2 -1446 13
rect -1428 -2 -1424 13
rect -1420 -2 -1416 13
rect -1412 18 -1408 33
rect -1381 17 -1377 33
rect -1393 13 -1388 17
rect -1381 13 -1373 17
rect -1412 -2 -1408 13
rect -1381 -2 -1377 13
rect -1614 -9 -1610 -6
rect -1595 -9 -1591 -6
rect -1554 -9 -1550 -6
rect -1532 -9 -1528 -6
rect -1458 -9 -1454 -6
rect -1436 -9 -1432 -6
rect -1389 -9 -1385 -6
rect -1614 -10 -1377 -9
rect -1614 -14 -1613 -10
rect -1609 -14 -1594 -10
rect -1590 -14 -1553 -10
rect -1549 -14 -1531 -10
rect -1527 -14 -1457 -10
rect -1453 -14 -1435 -10
rect -1431 -14 -1388 -10
rect -1384 -14 -1377 -10
rect -1614 -15 -1377 -14
rect -1600 -43 -1572 -39
rect -1568 -43 -1416 -39
rect -1624 -52 -1512 -48
rect -1508 -52 -1476 -48
rect -1382 -64 -1377 -15
rect -1733 -68 -1377 -64
rect -1733 -239 -1724 -68
rect -1626 -85 -1574 -81
rect -1570 -85 -1418 -81
rect -1626 -139 -1622 -85
rect -1602 -94 -1514 -90
rect -1510 -94 -1478 -90
rect -1354 -106 -1349 44
rect -1616 -107 -1349 -106
rect -1616 -111 -1615 -107
rect -1611 -111 -1596 -107
rect -1592 -111 -1555 -107
rect -1551 -111 -1533 -107
rect -1529 -111 -1459 -107
rect -1455 -111 -1437 -107
rect -1433 -111 -1390 -107
rect -1386 -111 -1349 -107
rect -1616 -112 -1349 -111
rect -1616 -115 -1612 -112
rect -1597 -115 -1593 -112
rect -1556 -115 -1552 -112
rect -1534 -115 -1530 -112
rect -1460 -115 -1456 -112
rect -1438 -115 -1434 -112
rect -1391 -115 -1387 -112
rect -1608 -138 -1604 -123
rect -1626 -143 -1615 -139
rect -1589 -139 -1585 -123
rect -1578 -139 -1574 -123
rect -1589 -143 -1574 -139
rect -1626 -204 -1622 -143
rect -1608 -158 -1604 -143
rect -1589 -158 -1585 -143
rect -1578 -158 -1574 -143
rect -1570 -138 -1566 -123
rect -1548 -139 -1544 -131
rect -1526 -139 -1522 -123
rect -1518 -139 -1514 -123
rect -1565 -143 -1555 -139
rect -1548 -143 -1541 -139
rect -1537 -143 -1533 -139
rect -1526 -143 -1514 -139
rect -1570 -158 -1566 -143
rect -1548 -154 -1544 -143
rect -1526 -158 -1522 -143
rect -1518 -158 -1514 -143
rect -1510 -138 -1506 -123
rect -1482 -138 -1478 -123
rect -1510 -158 -1506 -143
rect -1482 -158 -1478 -143
rect -1474 -139 -1470 -123
rect -1474 -143 -1466 -139
rect -1452 -139 -1448 -131
rect -1461 -143 -1459 -139
rect -1452 -143 -1445 -139
rect -1430 -139 -1426 -123
rect -1422 -139 -1418 -123
rect -1440 -143 -1437 -139
rect -1430 -143 -1418 -139
rect -1474 -158 -1470 -143
rect -1452 -154 -1448 -143
rect -1430 -158 -1426 -143
rect -1422 -158 -1418 -143
rect -1414 -138 -1410 -123
rect -1383 -139 -1379 -123
rect -1395 -143 -1390 -139
rect -1383 -143 -1375 -139
rect -1414 -158 -1410 -143
rect -1383 -158 -1379 -143
rect -1616 -165 -1612 -162
rect -1597 -165 -1593 -162
rect -1556 -165 -1552 -162
rect -1534 -165 -1530 -162
rect -1460 -165 -1456 -162
rect -1438 -165 -1434 -162
rect -1391 -165 -1387 -162
rect -1616 -166 -1379 -165
rect -1616 -170 -1615 -166
rect -1611 -170 -1596 -166
rect -1592 -170 -1555 -166
rect -1551 -170 -1533 -166
rect -1529 -170 -1459 -166
rect -1455 -170 -1437 -166
rect -1433 -170 -1390 -166
rect -1386 -170 -1379 -166
rect -1616 -171 -1379 -170
rect -1602 -199 -1574 -195
rect -1570 -199 -1418 -195
rect -1626 -208 -1514 -204
rect -1510 -208 -1478 -204
rect -1383 -239 -1379 -171
rect -1733 -243 -1379 -239
rect -1733 -452 -1724 -243
rect -1626 -293 -1574 -289
rect -1570 -293 -1418 -289
rect -1626 -347 -1622 -293
rect -1602 -302 -1514 -298
rect -1510 -302 -1478 -298
rect -1362 -314 -1358 -112
rect -1616 -315 -1358 -314
rect -1616 -319 -1615 -315
rect -1611 -319 -1596 -315
rect -1592 -319 -1555 -315
rect -1551 -319 -1533 -315
rect -1529 -319 -1459 -315
rect -1455 -319 -1437 -315
rect -1433 -319 -1390 -315
rect -1386 -319 -1358 -315
rect -1616 -320 -1358 -319
rect -1616 -323 -1612 -320
rect -1597 -323 -1593 -320
rect -1556 -323 -1552 -320
rect -1534 -323 -1530 -320
rect -1460 -323 -1456 -320
rect -1438 -323 -1434 -320
rect -1391 -323 -1387 -320
rect -1608 -346 -1604 -331
rect -1626 -351 -1615 -347
rect -1589 -347 -1585 -331
rect -1578 -347 -1574 -331
rect -1589 -351 -1574 -347
rect -1626 -412 -1622 -351
rect -1608 -366 -1604 -351
rect -1589 -366 -1585 -351
rect -1578 -366 -1574 -351
rect -1570 -346 -1566 -331
rect -1548 -347 -1544 -339
rect -1526 -347 -1522 -331
rect -1518 -347 -1514 -331
rect -1565 -351 -1555 -347
rect -1548 -351 -1541 -347
rect -1537 -351 -1533 -347
rect -1526 -351 -1514 -347
rect -1570 -366 -1566 -351
rect -1548 -362 -1544 -351
rect -1526 -366 -1522 -351
rect -1518 -366 -1514 -351
rect -1510 -346 -1506 -331
rect -1482 -346 -1478 -331
rect -1510 -366 -1506 -351
rect -1482 -366 -1478 -351
rect -1474 -347 -1470 -331
rect -1474 -351 -1466 -347
rect -1452 -347 -1448 -339
rect -1461 -351 -1459 -347
rect -1452 -351 -1445 -347
rect -1430 -347 -1426 -331
rect -1422 -347 -1418 -331
rect -1440 -351 -1437 -347
rect -1430 -351 -1418 -347
rect -1474 -366 -1470 -351
rect -1452 -362 -1448 -351
rect -1430 -366 -1426 -351
rect -1422 -366 -1418 -351
rect -1414 -346 -1410 -331
rect -1383 -347 -1379 -331
rect -1395 -351 -1390 -347
rect -1383 -351 -1375 -347
rect -1414 -366 -1410 -351
rect -1383 -366 -1379 -351
rect -1616 -373 -1612 -370
rect -1597 -373 -1593 -370
rect -1556 -373 -1552 -370
rect -1534 -373 -1530 -370
rect -1460 -373 -1456 -370
rect -1438 -373 -1434 -370
rect -1391 -373 -1387 -370
rect -1616 -374 -1379 -373
rect -1616 -378 -1615 -374
rect -1611 -378 -1596 -374
rect -1592 -378 -1555 -374
rect -1551 -378 -1533 -374
rect -1529 -378 -1459 -374
rect -1455 -378 -1437 -374
rect -1433 -378 -1390 -374
rect -1386 -378 -1379 -374
rect -1616 -379 -1379 -378
rect -1602 -407 -1574 -403
rect -1570 -407 -1418 -403
rect -1626 -416 -1514 -412
rect -1510 -416 -1478 -412
rect -1384 -452 -1379 -379
rect -1733 -457 -1379 -452
rect -1362 -390 -1358 -320
rect -861 -382 -857 -379
rect -853 -382 -849 -147
rect -517 -303 -513 9
rect -376 -138 -251 -134
rect -247 -138 53 -134
rect -441 -156 -52 -152
rect -445 -175 -441 -156
rect -437 -175 -433 -172
rect -364 -170 -317 -166
rect -364 -175 -360 -170
rect -392 -179 -364 -175
rect -351 -179 -348 -175
rect -321 -176 -317 -170
rect -235 -169 -188 -165
rect -235 -175 -231 -169
rect -263 -179 -235 -175
rect -222 -179 -219 -175
rect -192 -176 -188 -169
rect -56 -175 -52 -156
rect 49 -157 53 -138
rect 20 -161 145 -157
rect 149 -161 153 -157
rect -48 -175 -44 -172
rect 32 -171 79 -167
rect 32 -175 36 -171
rect 4 -179 32 -175
rect 45 -179 48 -175
rect 75 -176 79 -171
rect 161 -169 208 -165
rect 161 -175 165 -169
rect 133 -179 161 -175
rect 174 -179 177 -175
rect 204 -176 208 -169
rect 287 -183 292 106
rect -449 -184 292 -183
rect -449 -188 -441 -184
rect -437 -188 -384 -184
rect -380 -188 -325 -184
rect -321 -188 -308 -184
rect -304 -188 -255 -184
rect -251 -188 -196 -184
rect -192 -188 -179 -184
rect -175 -188 -143 -184
rect -139 -188 -118 -184
rect -114 -188 -52 -184
rect -48 -188 -35 -184
rect -31 -188 12 -184
rect 16 -188 71 -184
rect 75 -188 88 -184
rect 92 -188 141 -184
rect 145 -188 200 -184
rect 204 -188 217 -184
rect 221 -188 253 -184
rect 257 -188 278 -184
rect 282 -188 292 -184
rect -449 -189 292 -188
rect -449 -205 -445 -189
rect -433 -205 -429 -189
rect -400 -192 -396 -189
rect -384 -192 -380 -189
rect -360 -192 -356 -189
rect -441 -224 -437 -213
rect -441 -225 -429 -224
rect -441 -228 -399 -225
rect -433 -229 -399 -228
rect -392 -228 -388 -200
rect -376 -228 -372 -200
rect -364 -208 -352 -204
rect -348 -196 -336 -192
rect -326 -194 -322 -189
rect -308 -194 -304 -189
rect -299 -192 -295 -189
rect -271 -192 -267 -189
rect -255 -192 -251 -189
rect -231 -192 -227 -189
rect -344 -222 -340 -208
rect -352 -226 -332 -222
rect -433 -239 -429 -229
rect -449 -267 -445 -247
rect -392 -260 -388 -233
rect -376 -260 -372 -233
rect -352 -256 -348 -226
rect -317 -231 -313 -198
rect -291 -231 -287 -200
rect -272 -212 -270 -208
rect -263 -228 -259 -200
rect -247 -228 -243 -200
rect -235 -208 -223 -204
rect -219 -196 -207 -192
rect -197 -194 -193 -189
rect -179 -194 -175 -189
rect -170 -192 -166 -189
rect -144 -192 -140 -189
rect -118 -192 -114 -189
rect -215 -222 -211 -208
rect -223 -226 -203 -222
rect -317 -235 -298 -231
rect -291 -235 -284 -231
rect -307 -256 -303 -235
rect -400 -267 -396 -264
rect -384 -267 -380 -264
rect -368 -267 -364 -264
rect -336 -267 -332 -264
rect -291 -260 -287 -235
rect -263 -260 -259 -233
rect -247 -260 -243 -233
rect -223 -256 -219 -226
rect -188 -231 -184 -198
rect -162 -231 -158 -200
rect -127 -205 -123 -200
rect -108 -205 -104 -200
rect -135 -209 -116 -205
rect -108 -209 -73 -205
rect -188 -235 -169 -231
rect -162 -235 -142 -231
rect -178 -256 -174 -235
rect -327 -267 -323 -264
rect -299 -267 -295 -264
rect -271 -267 -267 -264
rect -255 -267 -251 -264
rect -239 -267 -235 -264
rect -207 -267 -203 -264
rect -162 -260 -158 -235
rect -135 -255 -131 -209
rect -108 -260 -104 -209
rect -60 -208 -56 -189
rect -44 -208 -40 -189
rect -36 -208 -32 -189
rect -4 -192 0 -189
rect 12 -192 16 -189
rect 36 -192 40 -189
rect -52 -227 -48 -216
rect -52 -230 -40 -227
rect -28 -228 -24 -216
rect 4 -228 8 -200
rect 20 -228 24 -200
rect 32 -208 44 -204
rect 48 -196 60 -192
rect 70 -194 74 -189
rect 88 -194 92 -189
rect 97 -192 101 -189
rect 125 -192 129 -189
rect 141 -192 145 -189
rect 165 -192 169 -189
rect 52 -222 56 -208
rect 44 -226 64 -222
rect -52 -231 -35 -230
rect -44 -234 -35 -231
rect -28 -232 -3 -228
rect -44 -242 -40 -234
rect -198 -267 -194 -264
rect -170 -267 -166 -264
rect -144 -267 -140 -263
rect -127 -267 -123 -263
rect -28 -246 -24 -232
rect -118 -267 -114 -264
rect -60 -267 -56 -250
rect -36 -267 -32 -250
rect 4 -260 8 -233
rect 20 -260 24 -233
rect 44 -256 48 -226
rect 79 -231 83 -198
rect 105 -231 109 -200
rect 124 -212 126 -208
rect 133 -228 137 -200
rect 149 -228 153 -200
rect 161 -208 173 -204
rect 177 -196 189 -192
rect 199 -194 203 -189
rect 217 -194 221 -189
rect 226 -192 230 -189
rect 252 -192 256 -189
rect 278 -192 282 -189
rect 181 -222 185 -208
rect 173 -226 193 -222
rect 79 -235 98 -231
rect 105 -235 112 -231
rect 89 -256 93 -235
rect -4 -267 0 -264
rect 12 -267 16 -264
rect 28 -267 32 -264
rect 60 -267 64 -264
rect 105 -260 109 -235
rect 133 -260 137 -233
rect 149 -260 153 -233
rect 173 -256 177 -226
rect 208 -231 212 -198
rect 234 -231 238 -200
rect 269 -205 273 -200
rect 288 -205 292 -200
rect 261 -209 280 -205
rect 288 -209 299 -205
rect 208 -235 227 -231
rect 234 -235 254 -231
rect 218 -256 222 -235
rect 69 -267 73 -264
rect 97 -267 101 -264
rect 125 -267 129 -264
rect 141 -267 145 -264
rect 157 -267 161 -264
rect 189 -267 193 -264
rect 234 -260 238 -235
rect 261 -255 265 -209
rect 288 -260 292 -209
rect 198 -267 202 -264
rect 226 -267 230 -264
rect 252 -267 256 -263
rect 269 -267 273 -263
rect 295 -263 299 -209
rect 278 -267 282 -264
rect -449 -268 292 -267
rect -449 -272 -448 -268
rect -444 -272 -399 -268
rect -395 -272 -326 -268
rect -322 -272 -308 -268
rect -304 -272 -298 -268
rect -294 -272 -270 -268
rect -266 -272 -197 -268
rect -193 -272 -179 -268
rect -175 -272 -169 -268
rect -165 -272 -136 -268
rect -132 -272 -118 -268
rect -114 -272 -59 -268
rect -55 -272 -35 -268
rect -31 -272 -3 -268
rect 1 -272 70 -268
rect 74 -272 88 -268
rect 92 -272 98 -268
rect 102 -272 126 -268
rect 130 -272 199 -268
rect 203 -272 217 -268
rect 221 -272 227 -268
rect 231 -272 260 -268
rect 264 -272 278 -268
rect 282 -272 292 -268
rect -449 -273 292 -272
rect -376 -281 -356 -277
rect -356 -288 -352 -281
rect -343 -281 -340 -277
rect -313 -288 -309 -280
rect -247 -281 -227 -277
rect -356 -292 -309 -288
rect -227 -288 -223 -281
rect -214 -281 -211 -277
rect -184 -288 -180 -280
rect -131 -282 -127 -280
rect 20 -281 40 -277
rect -227 -292 -180 -288
rect 40 -288 44 -281
rect 53 -281 56 -277
rect 83 -288 87 -280
rect 149 -281 169 -277
rect 40 -292 87 -288
rect 169 -288 173 -281
rect 182 -281 185 -277
rect 212 -288 216 -280
rect 265 -282 269 -280
rect 287 -280 292 -273
rect 287 -284 341 -280
rect 169 -292 216 -288
rect -517 -307 -439 -303
rect -773 -376 -726 -372
rect -773 -382 -769 -376
rect -801 -386 -773 -382
rect -760 -386 -757 -382
rect -730 -383 -726 -376
rect -644 -376 -597 -372
rect -644 -382 -640 -376
rect -672 -386 -644 -382
rect -631 -386 -628 -382
rect -601 -383 -597 -376
rect -451 -382 -447 -379
rect -443 -382 -439 -307
rect -423 -340 -419 -338
rect -103 -342 -99 -294
rect -246 -346 -99 -342
rect 28 -364 32 -360
rect -370 -376 -323 -372
rect -370 -382 -366 -376
rect -398 -386 -370 -382
rect -357 -386 -354 -382
rect -327 -383 -323 -376
rect -241 -376 -194 -372
rect -241 -382 -237 -376
rect -269 -386 -241 -382
rect -228 -386 -225 -382
rect -198 -383 -194 -376
rect -1362 -391 -110 -390
rect -1362 -395 -857 -391
rect -853 -395 -840 -391
rect -836 -395 -792 -391
rect -788 -395 -734 -391
rect -730 -395 -717 -391
rect -713 -395 -664 -391
rect -660 -395 -605 -391
rect -601 -395 -588 -391
rect -584 -395 -552 -391
rect -548 -395 -527 -391
rect -523 -395 -447 -391
rect -443 -395 -390 -391
rect -386 -395 -331 -391
rect -327 -395 -314 -391
rect -310 -395 -261 -391
rect -257 -395 -202 -391
rect -198 -395 -185 -391
rect -181 -395 -149 -391
rect -145 -395 -124 -391
rect -120 -395 -110 -391
rect -1733 -718 -1724 -457
rect -1629 -516 -1577 -512
rect -1573 -516 -1421 -512
rect -1629 -570 -1625 -516
rect -1605 -525 -1517 -521
rect -1513 -525 -1481 -521
rect -1362 -536 -1358 -395
rect -865 -396 -110 -395
rect -865 -415 -861 -396
rect -849 -415 -845 -396
rect -841 -415 -837 -396
rect -809 -399 -805 -396
rect -793 -399 -789 -396
rect -769 -399 -765 -396
rect -857 -434 -853 -423
rect -857 -437 -845 -434
rect -833 -435 -829 -423
rect -801 -435 -797 -407
rect -785 -435 -781 -407
rect -773 -415 -761 -411
rect -757 -403 -745 -399
rect -735 -401 -731 -396
rect -717 -401 -713 -396
rect -708 -399 -704 -396
rect -680 -399 -676 -396
rect -664 -399 -660 -396
rect -640 -399 -636 -396
rect -753 -429 -749 -415
rect -761 -433 -741 -429
rect -857 -438 -840 -437
rect -849 -441 -840 -438
rect -833 -439 -808 -435
rect -849 -449 -845 -441
rect -833 -453 -829 -439
rect -865 -474 -861 -457
rect -841 -474 -837 -457
rect -801 -467 -797 -440
rect -785 -467 -781 -440
rect -761 -463 -757 -433
rect -726 -438 -722 -405
rect -700 -438 -696 -407
rect -681 -419 -679 -415
rect -672 -435 -668 -407
rect -656 -435 -652 -407
rect -644 -415 -632 -411
rect -628 -403 -616 -399
rect -606 -401 -602 -396
rect -588 -401 -584 -396
rect -579 -399 -575 -396
rect -553 -399 -549 -396
rect -527 -399 -523 -396
rect -624 -429 -620 -415
rect -632 -433 -612 -429
rect -726 -442 -707 -438
rect -700 -442 -693 -438
rect -716 -463 -712 -442
rect -809 -474 -805 -471
rect -793 -474 -789 -471
rect -777 -474 -773 -471
rect -745 -474 -741 -471
rect -700 -467 -696 -442
rect -672 -467 -668 -440
rect -656 -467 -652 -440
rect -632 -463 -628 -433
rect -597 -438 -593 -405
rect -571 -438 -567 -407
rect -536 -412 -532 -407
rect -517 -412 -513 -407
rect -455 -412 -451 -396
rect -439 -412 -435 -396
rect -406 -399 -402 -396
rect -390 -399 -386 -396
rect -366 -399 -362 -396
rect -544 -416 -525 -412
rect -517 -416 -504 -412
rect -597 -442 -578 -438
rect -571 -442 -551 -438
rect -587 -463 -583 -442
rect -736 -474 -732 -471
rect -708 -474 -704 -471
rect -680 -474 -676 -471
rect -664 -474 -660 -471
rect -648 -474 -644 -471
rect -616 -474 -612 -471
rect -571 -467 -567 -442
rect -544 -462 -540 -416
rect -517 -467 -513 -416
rect -508 -451 -504 -416
rect -447 -431 -443 -420
rect -447 -432 -435 -431
rect -447 -435 -405 -432
rect -439 -436 -405 -435
rect -398 -435 -394 -407
rect -382 -435 -378 -407
rect -370 -415 -358 -411
rect -354 -403 -342 -399
rect -332 -401 -328 -396
rect -314 -401 -310 -396
rect -305 -399 -301 -396
rect -277 -399 -273 -396
rect -261 -399 -257 -396
rect -237 -399 -233 -396
rect -350 -429 -346 -415
rect -358 -433 -338 -429
rect -439 -446 -435 -436
rect -607 -474 -603 -471
rect -579 -474 -575 -471
rect -553 -474 -549 -470
rect -536 -474 -532 -470
rect -527 -474 -523 -471
rect -455 -474 -451 -454
rect -398 -467 -394 -440
rect -382 -467 -378 -440
rect -358 -463 -354 -433
rect -323 -438 -319 -405
rect -297 -438 -293 -407
rect -278 -419 -276 -415
rect -269 -435 -265 -407
rect -253 -435 -249 -407
rect -241 -415 -229 -411
rect -225 -403 -213 -399
rect -203 -401 -199 -396
rect -185 -401 -181 -396
rect -176 -399 -172 -396
rect -150 -399 -146 -396
rect -124 -399 -120 -396
rect -221 -429 -217 -415
rect -229 -433 -209 -429
rect -323 -442 -304 -438
rect -297 -442 -290 -438
rect -313 -463 -309 -442
rect -406 -474 -402 -471
rect -390 -474 -386 -471
rect -374 -474 -370 -471
rect -342 -474 -338 -471
rect -297 -467 -293 -442
rect -269 -467 -265 -440
rect -253 -467 -249 -440
rect -229 -463 -225 -433
rect -194 -438 -190 -405
rect -168 -438 -164 -407
rect -133 -412 -129 -407
rect -114 -412 -110 -407
rect -141 -416 -122 -412
rect -114 -416 -102 -412
rect -194 -442 -175 -438
rect -168 -442 -148 -438
rect -184 -463 -180 -442
rect -333 -474 -329 -471
rect -305 -474 -301 -471
rect -277 -474 -273 -471
rect -261 -474 -257 -471
rect -245 -474 -241 -471
rect -213 -474 -209 -471
rect -168 -467 -164 -442
rect -141 -462 -137 -416
rect -114 -467 -110 -416
rect -204 -474 -200 -471
rect -176 -474 -172 -471
rect -150 -474 -146 -470
rect -133 -474 -129 -470
rect -106 -464 -102 -416
rect -124 -474 -120 -471
rect 287 -474 292 -284
rect -865 -475 292 -474
rect -865 -479 -864 -475
rect -860 -479 -840 -475
rect -836 -479 -808 -475
rect -804 -479 -735 -475
rect -731 -479 -717 -475
rect -713 -479 -707 -475
rect -703 -479 -679 -475
rect -675 -479 -606 -475
rect -602 -479 -588 -475
rect -584 -479 -578 -475
rect -574 -479 -545 -475
rect -541 -479 -527 -475
rect -523 -479 -454 -475
rect -450 -479 -405 -475
rect -401 -479 -332 -475
rect -328 -479 -314 -475
rect -310 -479 -304 -475
rect -300 -479 -276 -475
rect -272 -479 -203 -475
rect -199 -479 -185 -475
rect -181 -479 -175 -475
rect -171 -479 -142 -475
rect -138 -479 -124 -475
rect -120 -479 292 -475
rect -865 -480 292 -479
rect -785 -488 -765 -484
rect -765 -495 -761 -488
rect -752 -488 -749 -484
rect -722 -495 -718 -487
rect -656 -488 -636 -484
rect -765 -499 -718 -495
rect -636 -495 -632 -488
rect -623 -488 -620 -484
rect -593 -495 -589 -487
rect -540 -489 -536 -487
rect -382 -488 -362 -484
rect -636 -499 -589 -495
rect -362 -495 -358 -488
rect -349 -488 -346 -484
rect -319 -495 -315 -487
rect -253 -488 -233 -484
rect -362 -499 -315 -495
rect -233 -495 -229 -488
rect -220 -488 -217 -484
rect -190 -495 -186 -487
rect -137 -489 -133 -487
rect -233 -499 -186 -495
rect -1362 -537 -1251 -536
rect -1619 -538 -1251 -537
rect -1619 -542 -1618 -538
rect -1614 -542 -1599 -538
rect -1595 -542 -1558 -538
rect -1554 -542 -1536 -538
rect -1532 -542 -1462 -538
rect -1458 -542 -1440 -538
rect -1436 -542 -1393 -538
rect -1389 -540 -1251 -538
rect -1389 -542 -1358 -540
rect -1619 -543 -1358 -542
rect -1619 -546 -1615 -543
rect -1600 -546 -1596 -543
rect -1559 -546 -1555 -543
rect -1537 -546 -1533 -543
rect -1463 -546 -1459 -543
rect -1441 -546 -1437 -543
rect -1394 -546 -1390 -543
rect -1611 -569 -1607 -554
rect -1629 -574 -1618 -570
rect -1592 -570 -1588 -554
rect -1581 -570 -1577 -554
rect -1592 -574 -1577 -570
rect -1629 -635 -1625 -574
rect -1611 -589 -1607 -574
rect -1592 -589 -1588 -574
rect -1581 -589 -1577 -574
rect -1573 -569 -1569 -554
rect -1551 -570 -1547 -562
rect -1529 -570 -1525 -554
rect -1521 -570 -1517 -554
rect -1568 -574 -1558 -570
rect -1551 -574 -1544 -570
rect -1540 -574 -1536 -570
rect -1529 -574 -1517 -570
rect -1573 -589 -1569 -574
rect -1551 -585 -1547 -574
rect -1529 -589 -1525 -574
rect -1521 -589 -1517 -574
rect -1513 -569 -1509 -554
rect -1485 -569 -1481 -554
rect -1513 -589 -1509 -574
rect -1485 -589 -1481 -574
rect -1477 -570 -1473 -554
rect -1477 -574 -1469 -570
rect -1455 -570 -1451 -562
rect -1464 -574 -1462 -570
rect -1455 -574 -1448 -570
rect -1433 -570 -1429 -554
rect -1425 -570 -1421 -554
rect -1443 -574 -1440 -570
rect -1433 -574 -1421 -570
rect -1477 -589 -1473 -574
rect -1455 -585 -1451 -574
rect -1433 -589 -1429 -574
rect -1425 -589 -1421 -574
rect -1417 -569 -1413 -554
rect -1386 -570 -1382 -554
rect -1398 -574 -1393 -570
rect -1386 -574 -1378 -570
rect -1417 -589 -1413 -574
rect -1386 -589 -1382 -574
rect -1619 -596 -1615 -593
rect -1600 -596 -1596 -593
rect -1559 -596 -1555 -593
rect -1537 -596 -1533 -593
rect -1463 -596 -1459 -593
rect -1441 -596 -1437 -593
rect -1394 -596 -1390 -593
rect -1619 -597 -1363 -596
rect -1619 -601 -1618 -597
rect -1614 -601 -1599 -597
rect -1595 -601 -1558 -597
rect -1554 -601 -1536 -597
rect -1532 -601 -1462 -597
rect -1458 -601 -1440 -597
rect -1436 -601 -1393 -597
rect -1389 -601 -1363 -597
rect -1619 -602 -1363 -601
rect -1605 -630 -1577 -626
rect -1573 -630 -1421 -626
rect -1629 -639 -1517 -635
rect -1513 -639 -1481 -635
rect -1367 -718 -1363 -602
rect -1255 -634 -1251 -540
rect -1214 -562 -1210 -558
rect -1085 -589 -543 -585
rect -1085 -600 -1081 -589
rect -1198 -620 -1151 -616
rect -1198 -626 -1194 -620
rect -1226 -630 -1198 -626
rect -1185 -630 -1182 -626
rect -1155 -627 -1151 -620
rect -1069 -620 -1022 -616
rect -1069 -626 -1065 -620
rect -1097 -630 -1069 -626
rect -1056 -630 -1053 -626
rect -1026 -627 -1022 -620
rect -850 -626 -846 -622
rect -818 -620 -771 -616
rect -818 -626 -814 -620
rect -846 -630 -818 -626
rect -805 -630 -802 -626
rect -775 -627 -771 -620
rect -689 -620 -642 -616
rect -689 -626 -685 -620
rect -717 -630 -689 -626
rect -676 -630 -673 -626
rect -646 -627 -642 -620
rect -1255 -635 -558 -634
rect -1255 -639 -1218 -635
rect -1214 -639 -1159 -635
rect -1155 -639 -1142 -635
rect -1138 -639 -1089 -635
rect -1085 -639 -1030 -635
rect -1026 -639 -1013 -635
rect -1009 -639 -977 -635
rect -973 -639 -952 -635
rect -948 -639 -838 -635
rect -834 -639 -779 -635
rect -775 -639 -762 -635
rect -758 -639 -709 -635
rect -705 -639 -650 -635
rect -646 -639 -633 -635
rect -629 -639 -597 -635
rect -593 -639 -572 -635
rect -568 -639 -558 -635
rect -1234 -640 -558 -639
rect -1234 -643 -1230 -640
rect -1218 -643 -1214 -640
rect -1194 -643 -1190 -640
rect -1250 -663 -1233 -659
rect -1226 -679 -1222 -651
rect -1210 -679 -1206 -651
rect -1198 -659 -1186 -655
rect -1182 -647 -1170 -643
rect -1160 -645 -1156 -640
rect -1142 -645 -1138 -640
rect -1133 -643 -1129 -640
rect -1105 -643 -1101 -640
rect -1089 -643 -1085 -640
rect -1065 -643 -1061 -640
rect -1178 -673 -1174 -659
rect -1186 -677 -1166 -673
rect -1226 -711 -1222 -684
rect -1210 -711 -1206 -684
rect -1186 -707 -1182 -677
rect -1151 -682 -1147 -649
rect -1125 -682 -1121 -651
rect -1106 -663 -1104 -659
rect -1097 -679 -1093 -651
rect -1081 -679 -1077 -651
rect -1069 -659 -1057 -655
rect -1053 -647 -1041 -643
rect -1031 -645 -1027 -640
rect -1013 -645 -1009 -640
rect -1004 -643 -1000 -640
rect -978 -643 -974 -640
rect -952 -643 -948 -640
rect -854 -643 -850 -640
rect -838 -643 -834 -640
rect -814 -643 -810 -640
rect -1049 -673 -1045 -659
rect -1057 -677 -1037 -673
rect -1151 -686 -1132 -682
rect -1125 -686 -1118 -682
rect -1141 -707 -1137 -686
rect -1234 -718 -1230 -715
rect -1218 -718 -1214 -715
rect -1202 -718 -1198 -715
rect -1170 -718 -1166 -715
rect -1125 -711 -1121 -686
rect -1097 -711 -1093 -684
rect -1081 -711 -1077 -684
rect -1057 -707 -1053 -677
rect -1022 -682 -1018 -649
rect -996 -682 -992 -651
rect -961 -656 -957 -651
rect -942 -656 -938 -651
rect -969 -660 -950 -656
rect -942 -660 -930 -656
rect -1022 -686 -1003 -682
rect -996 -686 -976 -682
rect -1012 -707 -1008 -686
rect -1161 -718 -1157 -715
rect -1133 -718 -1129 -715
rect -1105 -718 -1101 -715
rect -1089 -718 -1085 -715
rect -1073 -718 -1069 -715
rect -1041 -718 -1037 -715
rect -996 -711 -992 -686
rect -969 -706 -965 -660
rect -942 -711 -938 -660
rect -846 -679 -842 -651
rect -830 -679 -826 -651
rect -818 -659 -806 -655
rect -802 -647 -790 -643
rect -780 -645 -776 -640
rect -762 -645 -758 -640
rect -753 -643 -749 -640
rect -725 -643 -721 -640
rect -709 -643 -705 -640
rect -685 -643 -681 -640
rect -798 -673 -794 -659
rect -806 -677 -786 -673
rect -846 -711 -842 -684
rect -830 -711 -826 -684
rect -806 -707 -802 -677
rect -771 -682 -767 -649
rect -745 -682 -741 -651
rect -726 -663 -724 -659
rect -717 -679 -713 -651
rect -701 -679 -697 -651
rect -689 -659 -677 -655
rect -673 -647 -661 -643
rect -651 -645 -647 -640
rect -633 -645 -629 -640
rect -624 -643 -620 -640
rect -598 -643 -594 -640
rect -572 -643 -568 -640
rect -669 -673 -665 -659
rect -677 -677 -657 -673
rect -771 -686 -752 -682
rect -745 -686 -738 -682
rect -761 -707 -757 -686
rect -1032 -718 -1028 -715
rect -1004 -718 -1000 -715
rect -978 -718 -974 -714
rect -961 -718 -957 -714
rect -952 -718 -948 -715
rect -854 -718 -850 -715
rect -838 -718 -834 -715
rect -822 -718 -818 -715
rect -790 -718 -786 -715
rect -745 -711 -741 -686
rect -717 -711 -713 -684
rect -701 -711 -697 -684
rect -677 -707 -673 -677
rect -642 -682 -638 -649
rect -616 -682 -612 -651
rect -581 -656 -577 -651
rect -562 -656 -558 -651
rect -547 -656 -543 -589
rect -289 -604 -285 -600
rect -589 -660 -570 -656
rect -562 -660 -543 -656
rect -642 -686 -623 -682
rect -616 -686 -596 -682
rect -632 -707 -628 -686
rect -781 -718 -777 -715
rect -753 -718 -749 -715
rect -725 -718 -721 -715
rect -709 -718 -705 -715
rect -693 -718 -689 -715
rect -661 -718 -657 -715
rect -616 -711 -612 -686
rect -589 -706 -585 -660
rect -562 -711 -558 -660
rect -652 -718 -648 -715
rect -624 -718 -620 -715
rect -598 -718 -594 -714
rect -581 -718 -577 -714
rect -572 -718 -568 -715
rect 287 -718 292 -480
rect -1733 -719 292 -718
rect -1733 -723 -1233 -719
rect -1229 -723 -1160 -719
rect -1156 -723 -1142 -719
rect -1138 -723 -1132 -719
rect -1128 -723 -1104 -719
rect -1100 -723 -1031 -719
rect -1027 -723 -1013 -719
rect -1009 -723 -1003 -719
rect -999 -723 -970 -719
rect -966 -723 -952 -719
rect -948 -723 -853 -719
rect -849 -723 -780 -719
rect -776 -723 -762 -719
rect -758 -723 -752 -719
rect -748 -723 -724 -719
rect -720 -723 -651 -719
rect -647 -723 -633 -719
rect -629 -723 -623 -719
rect -619 -723 -590 -719
rect -586 -723 -572 -719
rect -568 -723 292 -719
rect -1733 -724 292 -723
rect -1733 -1191 -1724 -724
rect -1210 -732 -1190 -728
rect -1190 -739 -1186 -732
rect -1177 -732 -1174 -728
rect -1147 -739 -1143 -731
rect -1081 -732 -1061 -728
rect -1190 -743 -1143 -739
rect -1061 -739 -1057 -732
rect -1048 -732 -1045 -728
rect -1018 -739 -1014 -731
rect -965 -733 -961 -731
rect -830 -732 -810 -728
rect -1061 -743 -1014 -739
rect -810 -739 -806 -732
rect -797 -732 -794 -728
rect -767 -739 -763 -731
rect -701 -732 -681 -728
rect -810 -743 -763 -739
rect -681 -739 -677 -732
rect -668 -732 -665 -728
rect -638 -739 -634 -731
rect -585 -733 -581 -731
rect -681 -743 -634 -739
rect -1173 -816 -1169 -812
rect -783 -813 -780 -809
rect -272 -819 -268 -815
rect 358 -838 378 106
rect -967 -842 378 -838
rect -1210 -878 -1158 -874
rect -1154 -878 -1002 -874
rect -1210 -932 -1206 -878
rect -1186 -887 -1098 -883
rect -1094 -887 -1062 -883
rect -967 -899 -963 -842
rect -1200 -900 -963 -899
rect -1200 -904 -1199 -900
rect -1195 -904 -1181 -900
rect -1177 -904 -1139 -900
rect -1135 -904 -1117 -900
rect -1113 -904 -1043 -900
rect -1039 -904 -1021 -900
rect -1017 -904 -974 -900
rect -970 -904 -963 -900
rect -1200 -905 -963 -904
rect -820 -861 -768 -857
rect -764 -861 -612 -857
rect -1200 -908 -1196 -905
rect -1181 -908 -1177 -905
rect -1140 -908 -1136 -905
rect -1118 -908 -1114 -905
rect -1044 -908 -1040 -905
rect -1022 -908 -1018 -905
rect -975 -908 -971 -905
rect -1192 -931 -1188 -916
rect -1210 -936 -1199 -932
rect -1173 -932 -1169 -916
rect -1162 -932 -1158 -916
rect -1173 -936 -1158 -932
rect -1210 -997 -1206 -936
rect -1192 -951 -1188 -936
rect -1173 -951 -1169 -936
rect -1162 -951 -1158 -936
rect -1154 -931 -1150 -916
rect -1132 -932 -1128 -924
rect -1110 -932 -1106 -916
rect -1102 -932 -1098 -916
rect -1149 -936 -1139 -932
rect -1132 -936 -1125 -932
rect -1121 -936 -1117 -932
rect -1110 -936 -1098 -932
rect -1154 -951 -1150 -936
rect -1132 -947 -1128 -936
rect -1110 -951 -1106 -936
rect -1102 -951 -1098 -936
rect -1094 -931 -1090 -916
rect -1066 -931 -1062 -916
rect -1094 -951 -1090 -936
rect -1066 -951 -1062 -936
rect -1058 -932 -1054 -916
rect -1058 -936 -1050 -932
rect -1036 -932 -1032 -924
rect -1045 -936 -1043 -932
rect -1036 -936 -1029 -932
rect -1014 -932 -1010 -916
rect -1006 -932 -1002 -916
rect -1024 -936 -1021 -932
rect -1014 -936 -1002 -932
rect -1058 -951 -1054 -936
rect -1036 -947 -1032 -936
rect -1014 -951 -1010 -936
rect -1006 -951 -1002 -936
rect -998 -931 -994 -916
rect -967 -932 -963 -916
rect -820 -915 -816 -861
rect -796 -870 -708 -866
rect -704 -870 -672 -866
rect -577 -882 -573 -842
rect -810 -883 -573 -882
rect -810 -887 -809 -883
rect -805 -887 -791 -883
rect -787 -887 -749 -883
rect -745 -887 -727 -883
rect -723 -887 -653 -883
rect -649 -887 -631 -883
rect -627 -887 -584 -883
rect -580 -887 -573 -883
rect -810 -888 -573 -887
rect -328 -860 -276 -856
rect -272 -860 -120 -856
rect -810 -891 -806 -888
rect -791 -891 -787 -888
rect -750 -891 -746 -888
rect -728 -891 -724 -888
rect -654 -891 -650 -888
rect -632 -891 -628 -888
rect -585 -891 -581 -888
rect -802 -914 -798 -899
rect -820 -919 -809 -915
rect -783 -915 -779 -899
rect -772 -915 -768 -899
rect -783 -919 -768 -915
rect -979 -936 -974 -932
rect -967 -936 -938 -932
rect -998 -951 -994 -936
rect -967 -951 -963 -936
rect -1200 -958 -1196 -955
rect -1181 -958 -1177 -955
rect -1140 -958 -1136 -955
rect -1118 -958 -1114 -955
rect -1044 -958 -1040 -955
rect -1022 -958 -1018 -955
rect -975 -958 -971 -955
rect -1200 -959 -963 -958
rect -1200 -963 -1199 -959
rect -1195 -963 -1180 -959
rect -1176 -963 -1139 -959
rect -1135 -963 -1117 -959
rect -1113 -963 -1043 -959
rect -1039 -963 -1021 -959
rect -1017 -963 -974 -959
rect -970 -963 -963 -959
rect -1200 -964 -963 -963
rect -1186 -992 -1158 -988
rect -1154 -992 -1002 -988
rect -1210 -1001 -1098 -997
rect -1094 -1001 -1062 -997
rect -968 -1191 -963 -964
rect -820 -980 -816 -919
rect -802 -934 -798 -919
rect -783 -934 -779 -919
rect -772 -934 -768 -919
rect -764 -914 -760 -899
rect -742 -915 -738 -907
rect -720 -915 -716 -899
rect -712 -915 -708 -899
rect -759 -919 -749 -915
rect -742 -919 -735 -915
rect -731 -919 -727 -915
rect -720 -919 -708 -915
rect -764 -934 -760 -919
rect -742 -930 -738 -919
rect -720 -934 -716 -919
rect -712 -934 -708 -919
rect -704 -914 -700 -899
rect -676 -914 -672 -899
rect -704 -934 -700 -919
rect -676 -934 -672 -919
rect -668 -915 -664 -899
rect -668 -919 -660 -915
rect -646 -915 -642 -907
rect -655 -919 -653 -915
rect -646 -919 -639 -915
rect -624 -915 -620 -899
rect -616 -915 -612 -899
rect -634 -919 -631 -915
rect -624 -919 -612 -915
rect -668 -934 -664 -919
rect -646 -930 -642 -919
rect -624 -934 -620 -919
rect -616 -934 -612 -919
rect -608 -914 -604 -899
rect -577 -915 -573 -899
rect -328 -914 -324 -860
rect -304 -869 -216 -865
rect -212 -869 -180 -865
rect -85 -881 -81 -842
rect 120 -864 124 -860
rect -318 -882 -81 -881
rect -318 -886 -317 -882
rect -313 -886 -299 -882
rect -295 -886 -257 -882
rect -253 -886 -235 -882
rect -231 -886 -161 -882
rect -157 -886 -139 -882
rect -135 -886 -92 -882
rect -88 -886 -81 -882
rect -318 -887 -81 -886
rect 83 -875 135 -871
rect 139 -875 291 -871
rect -318 -890 -314 -887
rect -299 -890 -295 -887
rect -258 -890 -254 -887
rect -236 -890 -232 -887
rect -162 -890 -158 -887
rect -140 -890 -136 -887
rect -93 -890 -89 -887
rect -310 -913 -306 -898
rect -589 -919 -584 -915
rect -577 -919 -546 -915
rect -328 -918 -317 -914
rect -291 -914 -287 -898
rect -280 -914 -276 -898
rect -291 -918 -276 -914
rect -608 -934 -604 -919
rect -577 -934 -573 -919
rect -810 -941 -806 -938
rect -791 -941 -787 -938
rect -750 -941 -746 -938
rect -728 -941 -724 -938
rect -654 -941 -650 -938
rect -632 -941 -628 -938
rect -585 -941 -581 -938
rect -810 -942 -573 -941
rect -810 -946 -809 -942
rect -805 -946 -790 -942
rect -786 -946 -749 -942
rect -745 -946 -727 -942
rect -723 -946 -653 -942
rect -649 -946 -631 -942
rect -627 -946 -584 -942
rect -580 -946 -573 -942
rect -810 -947 -573 -946
rect -796 -975 -768 -971
rect -764 -975 -612 -971
rect -820 -984 -708 -980
rect -704 -984 -672 -980
rect -577 -1191 -573 -947
rect -328 -979 -324 -918
rect -310 -933 -306 -918
rect -291 -933 -287 -918
rect -280 -933 -276 -918
rect -272 -913 -268 -898
rect -250 -914 -246 -906
rect -228 -914 -224 -898
rect -220 -914 -216 -898
rect -267 -918 -257 -914
rect -250 -918 -243 -914
rect -239 -918 -235 -914
rect -228 -918 -216 -914
rect -272 -933 -268 -918
rect -250 -929 -246 -918
rect -228 -933 -224 -918
rect -220 -933 -216 -918
rect -212 -913 -208 -898
rect -184 -913 -180 -898
rect -212 -933 -208 -918
rect -184 -933 -180 -918
rect -176 -914 -172 -898
rect -176 -918 -168 -914
rect -154 -914 -150 -906
rect -163 -918 -161 -914
rect -154 -918 -147 -914
rect -132 -914 -128 -898
rect -124 -914 -120 -898
rect -142 -918 -139 -914
rect -132 -918 -120 -914
rect -176 -933 -172 -918
rect -154 -929 -150 -918
rect -132 -933 -128 -918
rect -124 -933 -120 -918
rect -116 -913 -112 -898
rect -85 -914 -81 -898
rect -97 -918 -92 -914
rect -85 -918 -77 -914
rect -116 -933 -112 -918
rect -85 -933 -81 -918
rect 83 -929 87 -875
rect 107 -884 195 -880
rect 199 -884 231 -880
rect 326 -896 330 -842
rect 93 -897 330 -896
rect 93 -901 94 -897
rect 98 -901 112 -897
rect 116 -901 154 -897
rect 158 -901 176 -897
rect 180 -901 250 -897
rect 254 -901 272 -897
rect 276 -901 319 -897
rect 323 -901 330 -897
rect 93 -902 330 -901
rect 93 -905 97 -902
rect 112 -905 116 -902
rect 153 -905 157 -902
rect 175 -905 179 -902
rect 249 -905 253 -902
rect 271 -905 275 -902
rect 318 -905 322 -902
rect 101 -928 105 -913
rect 83 -933 94 -929
rect 120 -929 124 -913
rect 131 -929 135 -913
rect 120 -933 135 -929
rect -318 -940 -314 -937
rect -299 -940 -295 -937
rect -258 -940 -254 -937
rect -236 -940 -232 -937
rect -162 -940 -158 -937
rect -140 -940 -136 -937
rect -93 -940 -89 -937
rect -318 -941 -81 -940
rect -318 -945 -317 -941
rect -313 -945 -298 -941
rect -294 -945 -257 -941
rect -253 -945 -235 -941
rect -231 -945 -161 -941
rect -157 -945 -139 -941
rect -135 -945 -92 -941
rect -88 -945 -81 -941
rect -318 -946 -81 -945
rect -304 -974 -276 -970
rect -272 -974 -120 -970
rect -328 -983 -216 -979
rect -212 -983 -180 -979
rect -86 -1191 -81 -946
rect 83 -994 87 -933
rect 101 -948 105 -933
rect 120 -948 124 -933
rect 131 -948 135 -933
rect 139 -928 143 -913
rect 161 -929 165 -921
rect 183 -929 187 -913
rect 191 -929 195 -913
rect 144 -933 154 -929
rect 161 -933 168 -929
rect 172 -933 176 -929
rect 183 -933 195 -929
rect 139 -948 143 -933
rect 161 -944 165 -933
rect 183 -948 187 -933
rect 191 -948 195 -933
rect 199 -928 203 -913
rect 227 -928 231 -913
rect 199 -948 203 -933
rect 227 -948 231 -933
rect 235 -929 239 -913
rect 235 -933 243 -929
rect 257 -929 261 -921
rect 248 -933 250 -929
rect 257 -933 264 -929
rect 279 -929 283 -913
rect 287 -929 291 -913
rect 269 -933 272 -929
rect 279 -933 291 -929
rect 235 -948 239 -933
rect 257 -944 261 -933
rect 279 -948 283 -933
rect 287 -948 291 -933
rect 295 -928 299 -913
rect 326 -929 330 -913
rect 314 -933 319 -929
rect 326 -933 334 -929
rect 295 -948 299 -933
rect 326 -948 330 -933
rect 93 -955 97 -952
rect 112 -955 116 -952
rect 153 -955 157 -952
rect 175 -955 179 -952
rect 249 -955 253 -952
rect 271 -955 275 -952
rect 318 -955 322 -952
rect 93 -956 330 -955
rect 93 -960 94 -956
rect 98 -960 113 -956
rect 117 -960 154 -956
rect 158 -960 176 -956
rect 180 -960 250 -956
rect 254 -960 272 -956
rect 276 -960 319 -956
rect 323 -960 330 -956
rect 93 -961 330 -960
rect 107 -989 135 -985
rect 139 -989 291 -985
rect 83 -998 195 -994
rect 199 -998 231 -994
rect 326 -1191 330 -961
rect 358 -1133 378 -842
rect -1733 -1201 397 -1191
<< metal2 >>
rect -1572 71 -1568 75
rect -1476 62 -1472 66
rect -1605 18 -1601 61
rect -1539 53 -1477 57
rect -1605 -38 -1601 13
rect -1539 17 -1535 53
rect -1481 18 -1477 53
rect -1443 53 -1394 57
rect -1443 18 -1439 53
rect -1398 18 -1394 53
rect -1369 13 -40 17
rect -1568 -9 -1564 13
rect -1507 -9 -1503 13
rect -1568 -13 -1503 -9
rect -1463 -16 -1459 13
rect -1411 -16 -1407 13
rect -1463 -20 -1407 -16
rect -1572 -43 -1568 -39
rect -1416 -43 -1412 -39
rect -1476 -52 -1472 -48
rect -1624 -58 -1620 -56
rect -1645 -62 -1620 -58
rect -1645 -216 -1639 -62
rect -1574 -85 -1570 -81
rect -1478 -94 -1474 -90
rect -1607 -138 -1603 -95
rect -1541 -103 -1479 -99
rect -1607 -194 -1603 -143
rect -1541 -139 -1537 -103
rect -1483 -138 -1479 -103
rect -1445 -103 -1396 -99
rect -1445 -138 -1441 -103
rect -1400 -138 -1396 -103
rect -1371 -143 -433 -139
rect -1570 -165 -1566 -143
rect -1509 -165 -1505 -143
rect -1570 -169 -1505 -165
rect -1465 -172 -1461 -143
rect -1413 -172 -1409 -143
rect -1465 -176 -1409 -172
rect -1341 -156 -445 -152
rect -1574 -199 -1570 -195
rect -1418 -199 -1414 -195
rect -1478 -208 -1474 -204
rect -1626 -216 -1622 -212
rect -1645 -220 -1622 -216
rect -1645 -425 -1639 -220
rect -1574 -293 -1570 -289
rect -1478 -302 -1474 -298
rect -1607 -346 -1603 -303
rect -1541 -311 -1479 -307
rect -1607 -402 -1603 -351
rect -1541 -347 -1537 -311
rect -1483 -346 -1479 -311
rect -1445 -311 -1396 -307
rect -1445 -346 -1441 -311
rect -1400 -346 -1396 -311
rect -1341 -347 -1337 -156
rect -437 -168 -433 -143
rect -48 -168 -44 13
rect 157 -161 340 -157
rect -355 -183 -351 -179
rect -226 -183 -222 -179
rect 41 -183 45 -179
rect 170 -183 174 -179
rect -375 -187 -351 -183
rect -246 -187 -222 -183
rect 21 -187 45 -183
rect 150 -187 174 -183
rect -375 -228 -371 -187
rect -277 -223 -273 -213
rect -327 -227 -273 -223
rect -246 -228 -242 -187
rect -198 -227 -99 -223
rect -391 -269 -387 -233
rect -391 -273 -344 -269
rect -348 -277 -344 -273
rect -283 -294 -279 -236
rect -262 -269 -258 -233
rect -262 -273 -215 -269
rect -219 -277 -215 -273
rect -132 -294 -128 -287
rect -103 -290 -99 -227
rect -283 -298 -128 -294
rect -77 -305 -73 -213
rect 21 -228 25 -187
rect 119 -223 123 -213
rect 69 -227 123 -223
rect 150 -228 154 -187
rect 198 -227 329 -223
rect 5 -269 9 -233
rect 5 -273 52 -269
rect 48 -277 52 -273
rect 113 -294 117 -236
rect 134 -269 138 -233
rect 134 -273 181 -269
rect 177 -277 181 -273
rect 264 -294 268 -287
rect 113 -298 268 -294
rect -423 -309 -73 -305
rect -1371 -351 -1337 -347
rect -1295 -323 -446 -319
rect -1570 -373 -1566 -351
rect -1509 -373 -1505 -351
rect -1570 -377 -1505 -373
rect -1465 -380 -1461 -351
rect -1413 -380 -1409 -351
rect -1465 -384 -1409 -380
rect -1574 -407 -1570 -403
rect -1418 -407 -1414 -403
rect -1478 -416 -1474 -412
rect -1626 -425 -1622 -420
rect -1645 -429 -1622 -425
rect -1645 -650 -1639 -429
rect -1577 -516 -1573 -512
rect -1481 -525 -1477 -521
rect -1610 -569 -1606 -526
rect -1544 -534 -1482 -530
rect -1610 -625 -1606 -574
rect -1544 -570 -1540 -534
rect -1486 -569 -1482 -534
rect -1448 -534 -1399 -530
rect -1448 -569 -1444 -534
rect -1403 -569 -1399 -534
rect -1295 -570 -1291 -323
rect -861 -375 -857 -323
rect -451 -375 -447 -323
rect -423 -334 -419 -309
rect 295 -360 299 -267
rect 36 -364 299 -360
rect -764 -390 -760 -386
rect -635 -390 -631 -386
rect -361 -390 -357 -386
rect -232 -390 -228 -386
rect -784 -394 -760 -390
rect -655 -394 -631 -390
rect -381 -394 -357 -390
rect -252 -394 -228 -390
rect -784 -435 -780 -394
rect -686 -430 -682 -420
rect -736 -434 -682 -430
rect -655 -435 -651 -394
rect -607 -434 -468 -430
rect -800 -476 -796 -440
rect -800 -480 -753 -476
rect -757 -484 -753 -480
rect -692 -501 -688 -443
rect -671 -476 -667 -440
rect -671 -480 -624 -476
rect -628 -484 -624 -480
rect -541 -501 -537 -494
rect -692 -505 -537 -501
rect -508 -515 -504 -455
rect -1214 -519 -504 -515
rect -1214 -554 -1210 -519
rect -473 -538 -468 -434
rect -381 -435 -377 -394
rect -283 -430 -279 -420
rect -333 -434 -279 -430
rect -252 -435 -248 -394
rect -204 -434 -83 -430
rect -397 -476 -393 -440
rect -397 -480 -350 -476
rect -354 -484 -350 -480
rect -289 -501 -285 -443
rect -268 -476 -264 -440
rect -268 -480 -221 -476
rect -225 -484 -221 -480
rect -138 -501 -134 -494
rect -289 -505 -134 -501
rect -850 -542 -468 -538
rect -1374 -574 -1291 -570
rect -1573 -596 -1569 -574
rect -1512 -596 -1508 -574
rect -1573 -600 -1508 -596
rect -1468 -603 -1464 -574
rect -1416 -603 -1412 -574
rect -1468 -607 -1412 -603
rect -850 -618 -846 -542
rect -106 -600 -102 -468
rect -281 -604 -102 -600
rect -1577 -630 -1573 -626
rect -1421 -630 -1417 -626
rect -1189 -634 -1185 -630
rect -1060 -634 -1056 -630
rect -809 -634 -805 -630
rect -680 -634 -676 -630
rect -1481 -639 -1477 -635
rect -1209 -638 -1185 -634
rect -1080 -638 -1056 -634
rect -829 -638 -805 -634
rect -700 -638 -676 -634
rect -1626 -650 -1622 -643
rect -1645 -654 -1622 -650
rect -1645 -1015 -1639 -654
rect -1209 -679 -1205 -638
rect -1111 -674 -1107 -664
rect -1161 -678 -1107 -674
rect -1080 -679 -1076 -638
rect -1032 -678 -922 -674
rect -1225 -720 -1221 -684
rect -1225 -724 -1178 -720
rect -1182 -728 -1178 -724
rect -1117 -745 -1113 -687
rect -1096 -720 -1092 -684
rect -1096 -724 -1049 -720
rect -1053 -728 -1049 -724
rect -966 -745 -962 -738
rect -1117 -749 -962 -745
rect -926 -812 -922 -678
rect -829 -679 -825 -638
rect -731 -674 -727 -664
rect -781 -678 -727 -674
rect -700 -679 -696 -638
rect -652 -678 -543 -674
rect -845 -720 -841 -684
rect -845 -724 -798 -720
rect -802 -728 -798 -724
rect -737 -737 -733 -687
rect -716 -720 -712 -684
rect -716 -724 -669 -720
rect -673 -728 -669 -724
rect -737 -738 -586 -737
rect -737 -741 -582 -738
rect -737 -743 -733 -741
rect -586 -743 -582 -741
rect -547 -809 -543 -678
rect -1165 -816 -922 -812
rect -776 -813 -543 -809
rect -87 -815 -83 -434
rect 325 -749 329 -227
rect 336 -276 340 -161
rect -264 -819 -83 -815
rect 270 -753 329 -749
rect -768 -861 -764 -857
rect -276 -860 -272 -856
rect 270 -860 274 -753
rect 128 -864 274 -860
rect -672 -870 -668 -866
rect -180 -869 -176 -865
rect -1158 -878 -1154 -874
rect -1062 -887 -1058 -883
rect -1191 -931 -1187 -888
rect -1125 -896 -1063 -892
rect -1191 -987 -1187 -936
rect -1125 -932 -1121 -896
rect -1067 -931 -1063 -896
rect -1029 -896 -980 -892
rect -1029 -931 -1025 -896
rect -984 -931 -980 -896
rect -801 -914 -797 -871
rect -735 -879 -673 -875
rect -1154 -958 -1150 -936
rect -1093 -958 -1089 -936
rect -1154 -962 -1089 -958
rect -1049 -965 -1045 -936
rect -997 -965 -993 -936
rect -1049 -969 -993 -965
rect -801 -970 -797 -919
rect -735 -915 -731 -879
rect -677 -914 -673 -879
rect -639 -879 -590 -875
rect -639 -914 -635 -879
rect -594 -914 -590 -879
rect -309 -913 -305 -870
rect -243 -878 -181 -874
rect -764 -941 -760 -919
rect -703 -941 -699 -919
rect -764 -945 -699 -941
rect -659 -948 -655 -919
rect -607 -948 -603 -919
rect -659 -952 -603 -948
rect -309 -969 -305 -918
rect -243 -914 -239 -878
rect -185 -913 -181 -878
rect -147 -878 -98 -874
rect 135 -875 139 -871
rect -147 -913 -143 -878
rect -102 -913 -98 -878
rect 231 -884 235 -880
rect -272 -940 -268 -918
rect -211 -940 -207 -918
rect -272 -944 -207 -940
rect -167 -947 -163 -918
rect -115 -947 -111 -918
rect 102 -928 106 -885
rect 168 -893 230 -889
rect -167 -951 -111 -947
rect -768 -975 -764 -971
rect -612 -975 -608 -971
rect -276 -974 -272 -970
rect -120 -974 -116 -970
rect -672 -984 -668 -980
rect -180 -983 -176 -979
rect -1158 -992 -1154 -988
rect -1002 -992 -998 -988
rect -1062 -1001 -1058 -997
rect -1210 -1015 -1206 -1006
rect -811 -1015 -807 -988
rect -323 -1015 -319 -987
rect 102 -984 106 -933
rect 168 -929 172 -893
rect 226 -928 230 -893
rect 264 -893 313 -889
rect 264 -928 268 -893
rect 309 -928 313 -893
rect 139 -955 143 -933
rect 200 -955 204 -933
rect 139 -959 204 -955
rect 244 -962 248 -933
rect 296 -962 300 -933
rect 244 -966 300 -962
rect 135 -989 139 -985
rect 291 -989 295 -985
rect 231 -998 235 -994
rect 87 -1015 91 -1002
rect -1645 -1019 91 -1015
<< ntransistor >>
rect -1609 -6 -1607 -2
rect -1590 -6 -1588 -2
rect -1571 -6 -1569 -2
rect -1549 -6 -1547 2
rect -1527 -6 -1525 -2
rect -1511 -6 -1509 -2
rect -1475 -6 -1473 -2
rect -1453 -6 -1451 2
rect -1431 -6 -1429 -2
rect -1415 -6 -1413 -2
rect -1384 -6 -1382 -2
rect -1611 -162 -1609 -158
rect -1592 -162 -1590 -158
rect -1573 -162 -1571 -158
rect -1551 -162 -1549 -154
rect -1529 -162 -1527 -158
rect -1513 -162 -1511 -158
rect -1477 -162 -1475 -158
rect -1455 -162 -1453 -154
rect -1433 -162 -1431 -158
rect -1417 -162 -1415 -158
rect -1386 -162 -1384 -158
rect -444 -247 -442 -239
rect -436 -247 -434 -239
rect -395 -264 -393 -260
rect -379 -264 -377 -260
rect -363 -264 -361 -256
rect -355 -264 -353 -256
rect -347 -264 -345 -256
rect -339 -264 -337 -256
rect -320 -264 -318 -256
rect -312 -264 -310 -256
rect -294 -264 -292 -260
rect -266 -264 -264 -260
rect -250 -264 -248 -260
rect -234 -264 -232 -256
rect -226 -264 -224 -256
rect -218 -264 -216 -256
rect -210 -264 -208 -256
rect -191 -264 -189 -256
rect -183 -264 -181 -256
rect -165 -264 -163 -260
rect -138 -263 -136 -255
rect -130 -263 -128 -255
rect -55 -250 -53 -242
rect -47 -250 -45 -242
rect -31 -250 -29 -246
rect -112 -264 -110 -260
rect 1 -264 3 -260
rect 17 -264 19 -260
rect 33 -264 35 -256
rect 41 -264 43 -256
rect 49 -264 51 -256
rect 57 -264 59 -256
rect 76 -264 78 -256
rect 84 -264 86 -256
rect 102 -264 104 -260
rect 130 -264 132 -260
rect 146 -264 148 -260
rect 162 -264 164 -256
rect 170 -264 172 -256
rect 178 -264 180 -256
rect 186 -264 188 -256
rect 205 -264 207 -256
rect 213 -264 215 -256
rect 231 -264 233 -260
rect 258 -263 260 -255
rect 266 -263 268 -255
rect 284 -264 286 -260
rect -1611 -370 -1609 -366
rect -1592 -370 -1590 -366
rect -1573 -370 -1571 -366
rect -1551 -370 -1549 -362
rect -1529 -370 -1527 -366
rect -1513 -370 -1511 -366
rect -1477 -370 -1475 -366
rect -1455 -370 -1453 -362
rect -1433 -370 -1431 -366
rect -1417 -370 -1415 -366
rect -1386 -370 -1384 -366
rect -860 -457 -858 -449
rect -852 -457 -850 -449
rect -836 -457 -834 -453
rect -804 -471 -802 -467
rect -788 -471 -786 -467
rect -772 -471 -770 -463
rect -764 -471 -762 -463
rect -756 -471 -754 -463
rect -748 -471 -746 -463
rect -729 -471 -727 -463
rect -721 -471 -719 -463
rect -703 -471 -701 -467
rect -675 -471 -673 -467
rect -659 -471 -657 -467
rect -643 -471 -641 -463
rect -635 -471 -633 -463
rect -627 -471 -625 -463
rect -619 -471 -617 -463
rect -600 -471 -598 -463
rect -592 -471 -590 -463
rect -574 -471 -572 -467
rect -547 -470 -545 -462
rect -539 -470 -537 -462
rect -450 -454 -448 -446
rect -442 -454 -440 -446
rect -521 -471 -519 -467
rect -401 -471 -399 -467
rect -385 -471 -383 -467
rect -369 -471 -367 -463
rect -361 -471 -359 -463
rect -353 -471 -351 -463
rect -345 -471 -343 -463
rect -326 -471 -324 -463
rect -318 -471 -316 -463
rect -300 -471 -298 -467
rect -272 -471 -270 -467
rect -256 -471 -254 -467
rect -240 -471 -238 -463
rect -232 -471 -230 -463
rect -224 -471 -222 -463
rect -216 -471 -214 -463
rect -197 -471 -195 -463
rect -189 -471 -187 -463
rect -171 -471 -169 -467
rect -144 -470 -142 -462
rect -136 -470 -134 -462
rect -118 -471 -116 -467
rect -1614 -593 -1612 -589
rect -1595 -593 -1593 -589
rect -1576 -593 -1574 -589
rect -1554 -593 -1552 -585
rect -1532 -593 -1530 -589
rect -1516 -593 -1514 -589
rect -1480 -593 -1478 -589
rect -1458 -593 -1456 -585
rect -1436 -593 -1434 -589
rect -1420 -593 -1418 -589
rect -1389 -593 -1387 -589
rect -1229 -715 -1227 -711
rect -1213 -715 -1211 -711
rect -1197 -715 -1195 -707
rect -1189 -715 -1187 -707
rect -1181 -715 -1179 -707
rect -1173 -715 -1171 -707
rect -1154 -715 -1152 -707
rect -1146 -715 -1144 -707
rect -1128 -715 -1126 -711
rect -1100 -715 -1098 -711
rect -1084 -715 -1082 -711
rect -1068 -715 -1066 -707
rect -1060 -715 -1058 -707
rect -1052 -715 -1050 -707
rect -1044 -715 -1042 -707
rect -1025 -715 -1023 -707
rect -1017 -715 -1015 -707
rect -999 -715 -997 -711
rect -972 -714 -970 -706
rect -964 -714 -962 -706
rect -946 -715 -944 -711
rect -849 -715 -847 -711
rect -833 -715 -831 -711
rect -817 -715 -815 -707
rect -809 -715 -807 -707
rect -801 -715 -799 -707
rect -793 -715 -791 -707
rect -774 -715 -772 -707
rect -766 -715 -764 -707
rect -748 -715 -746 -711
rect -720 -715 -718 -711
rect -704 -715 -702 -711
rect -688 -715 -686 -707
rect -680 -715 -678 -707
rect -672 -715 -670 -707
rect -664 -715 -662 -707
rect -645 -715 -643 -707
rect -637 -715 -635 -707
rect -619 -715 -617 -711
rect -592 -714 -590 -706
rect -584 -714 -582 -706
rect -566 -715 -564 -711
rect -1195 -955 -1193 -951
rect -1176 -955 -1174 -951
rect -1157 -955 -1155 -951
rect -1135 -955 -1133 -947
rect -1113 -955 -1111 -951
rect -1097 -955 -1095 -951
rect -1061 -955 -1059 -951
rect -1039 -955 -1037 -947
rect -805 -938 -803 -934
rect -786 -938 -784 -934
rect -767 -938 -765 -934
rect -745 -938 -743 -930
rect -723 -938 -721 -934
rect -707 -938 -705 -934
rect -671 -938 -669 -934
rect -649 -938 -647 -930
rect -627 -938 -625 -934
rect -611 -938 -609 -934
rect -580 -938 -578 -934
rect -313 -937 -311 -933
rect -294 -937 -292 -933
rect -275 -937 -273 -933
rect -253 -937 -251 -929
rect -231 -937 -229 -933
rect -215 -937 -213 -933
rect -179 -937 -177 -933
rect -157 -937 -155 -929
rect -135 -937 -133 -933
rect -119 -937 -117 -933
rect -88 -937 -86 -933
rect -1017 -955 -1015 -951
rect -1001 -955 -999 -951
rect -970 -955 -968 -951
rect 98 -952 100 -948
rect 117 -952 119 -948
rect 136 -952 138 -948
rect 158 -952 160 -944
rect 180 -952 182 -948
rect 196 -952 198 -948
rect 232 -952 234 -948
rect 254 -952 256 -944
rect 276 -952 278 -948
rect 292 -952 294 -948
rect 323 -952 325 -948
<< ptransistor >>
rect -1609 33 -1607 41
rect -1590 33 -1588 41
rect -1571 33 -1569 41
rect -1549 25 -1547 41
rect -1527 33 -1525 41
rect -1511 33 -1509 41
rect -1475 33 -1473 41
rect -1453 25 -1451 41
rect -1431 33 -1429 41
rect -1415 33 -1413 41
rect -1384 33 -1382 41
rect -1611 -123 -1609 -115
rect -1592 -123 -1590 -115
rect -1573 -123 -1571 -115
rect -1551 -131 -1549 -115
rect -1529 -123 -1527 -115
rect -1513 -123 -1511 -115
rect -1477 -123 -1475 -115
rect -1455 -131 -1453 -115
rect -1433 -123 -1431 -115
rect -1417 -123 -1415 -115
rect -1386 -123 -1384 -115
rect -395 -200 -393 -192
rect -379 -200 -377 -192
rect -444 -213 -442 -205
rect -436 -213 -434 -205
rect -363 -208 -361 -192
rect -355 -208 -353 -192
rect -347 -208 -345 -192
rect -339 -208 -337 -192
rect -320 -200 -318 -192
rect -312 -200 -310 -192
rect -294 -200 -292 -192
rect -266 -200 -264 -192
rect -250 -200 -248 -192
rect -234 -208 -232 -192
rect -226 -208 -224 -192
rect -218 -208 -216 -192
rect -210 -208 -208 -192
rect -191 -200 -189 -192
rect -183 -200 -181 -192
rect -165 -200 -163 -192
rect -138 -200 -136 -192
rect -130 -200 -128 -192
rect -112 -200 -110 -192
rect 1 -200 3 -192
rect 17 -200 19 -192
rect -55 -216 -53 -208
rect -47 -216 -45 -208
rect -31 -216 -29 -208
rect 33 -208 35 -192
rect 41 -208 43 -192
rect 49 -208 51 -192
rect 57 -208 59 -192
rect 76 -200 78 -192
rect 84 -200 86 -192
rect 102 -200 104 -192
rect 130 -200 132 -192
rect 146 -200 148 -192
rect 162 -208 164 -192
rect 170 -208 172 -192
rect 178 -208 180 -192
rect 186 -208 188 -192
rect 205 -200 207 -192
rect 213 -200 215 -192
rect 231 -200 233 -192
rect 258 -200 260 -192
rect 266 -200 268 -192
rect 284 -200 286 -192
rect -1611 -331 -1609 -323
rect -1592 -331 -1590 -323
rect -1573 -331 -1571 -323
rect -1551 -339 -1549 -323
rect -1529 -331 -1527 -323
rect -1513 -331 -1511 -323
rect -1477 -331 -1475 -323
rect -1455 -339 -1453 -323
rect -1433 -331 -1431 -323
rect -1417 -331 -1415 -323
rect -1386 -331 -1384 -323
rect -804 -407 -802 -399
rect -788 -407 -786 -399
rect -860 -423 -858 -415
rect -852 -423 -850 -415
rect -836 -423 -834 -415
rect -772 -415 -770 -399
rect -764 -415 -762 -399
rect -756 -415 -754 -399
rect -748 -415 -746 -399
rect -729 -407 -727 -399
rect -721 -407 -719 -399
rect -703 -407 -701 -399
rect -675 -407 -673 -399
rect -659 -407 -657 -399
rect -643 -415 -641 -399
rect -635 -415 -633 -399
rect -627 -415 -625 -399
rect -619 -415 -617 -399
rect -600 -407 -598 -399
rect -592 -407 -590 -399
rect -574 -407 -572 -399
rect -547 -407 -545 -399
rect -539 -407 -537 -399
rect -521 -407 -519 -399
rect -401 -407 -399 -399
rect -385 -407 -383 -399
rect -450 -420 -448 -412
rect -442 -420 -440 -412
rect -369 -415 -367 -399
rect -361 -415 -359 -399
rect -353 -415 -351 -399
rect -345 -415 -343 -399
rect -326 -407 -324 -399
rect -318 -407 -316 -399
rect -300 -407 -298 -399
rect -272 -407 -270 -399
rect -256 -407 -254 -399
rect -240 -415 -238 -399
rect -232 -415 -230 -399
rect -224 -415 -222 -399
rect -216 -415 -214 -399
rect -197 -407 -195 -399
rect -189 -407 -187 -399
rect -171 -407 -169 -399
rect -144 -407 -142 -399
rect -136 -407 -134 -399
rect -118 -407 -116 -399
rect -1614 -554 -1612 -546
rect -1595 -554 -1593 -546
rect -1576 -554 -1574 -546
rect -1554 -562 -1552 -546
rect -1532 -554 -1530 -546
rect -1516 -554 -1514 -546
rect -1480 -554 -1478 -546
rect -1458 -562 -1456 -546
rect -1436 -554 -1434 -546
rect -1420 -554 -1418 -546
rect -1389 -554 -1387 -546
rect -1229 -651 -1227 -643
rect -1213 -651 -1211 -643
rect -1197 -659 -1195 -643
rect -1189 -659 -1187 -643
rect -1181 -659 -1179 -643
rect -1173 -659 -1171 -643
rect -1154 -651 -1152 -643
rect -1146 -651 -1144 -643
rect -1128 -651 -1126 -643
rect -1100 -651 -1098 -643
rect -1084 -651 -1082 -643
rect -1068 -659 -1066 -643
rect -1060 -659 -1058 -643
rect -1052 -659 -1050 -643
rect -1044 -659 -1042 -643
rect -1025 -651 -1023 -643
rect -1017 -651 -1015 -643
rect -999 -651 -997 -643
rect -972 -651 -970 -643
rect -964 -651 -962 -643
rect -946 -651 -944 -643
rect -849 -651 -847 -643
rect -833 -651 -831 -643
rect -817 -659 -815 -643
rect -809 -659 -807 -643
rect -801 -659 -799 -643
rect -793 -659 -791 -643
rect -774 -651 -772 -643
rect -766 -651 -764 -643
rect -748 -651 -746 -643
rect -720 -651 -718 -643
rect -704 -651 -702 -643
rect -688 -659 -686 -643
rect -680 -659 -678 -643
rect -672 -659 -670 -643
rect -664 -659 -662 -643
rect -645 -651 -643 -643
rect -637 -651 -635 -643
rect -619 -651 -617 -643
rect -592 -651 -590 -643
rect -584 -651 -582 -643
rect -566 -651 -564 -643
rect -805 -899 -803 -891
rect -786 -899 -784 -891
rect -767 -899 -765 -891
rect -1195 -916 -1193 -908
rect -1176 -916 -1174 -908
rect -1157 -916 -1155 -908
rect -1135 -924 -1133 -908
rect -1113 -916 -1111 -908
rect -1097 -916 -1095 -908
rect -1061 -916 -1059 -908
rect -1039 -924 -1037 -908
rect -1017 -916 -1015 -908
rect -1001 -916 -999 -908
rect -970 -916 -968 -908
rect -745 -907 -743 -891
rect -723 -899 -721 -891
rect -707 -899 -705 -891
rect -671 -899 -669 -891
rect -649 -907 -647 -891
rect -627 -899 -625 -891
rect -611 -899 -609 -891
rect -580 -899 -578 -891
rect -313 -898 -311 -890
rect -294 -898 -292 -890
rect -275 -898 -273 -890
rect -253 -906 -251 -890
rect -231 -898 -229 -890
rect -215 -898 -213 -890
rect -179 -898 -177 -890
rect -157 -906 -155 -890
rect -135 -898 -133 -890
rect -119 -898 -117 -890
rect -88 -898 -86 -890
rect 98 -913 100 -905
rect 117 -913 119 -905
rect 136 -913 138 -905
rect 158 -921 160 -905
rect 180 -913 182 -905
rect 196 -913 198 -905
rect 232 -913 234 -905
rect 254 -921 256 -905
rect 276 -913 278 -905
rect 292 -913 294 -905
rect 323 -913 325 -905
<< polycontact >>
rect -1572 71 -1568 75
rect -1416 71 -1412 75
rect -1512 62 -1508 66
rect -1476 62 -1472 66
rect -1613 13 -1609 17
rect -1594 13 -1590 17
rect -1553 13 -1549 17
rect -1531 13 -1527 17
rect -1457 13 -1453 17
rect -1435 13 -1431 17
rect -1388 13 -1384 17
rect -1572 -43 -1568 -39
rect -1416 -43 -1412 -39
rect -1512 -52 -1508 -48
rect -1476 -52 -1472 -48
rect -1574 -85 -1570 -81
rect -1418 -85 -1414 -81
rect -1514 -94 -1510 -90
rect -1478 -94 -1474 -90
rect -1615 -143 -1611 -139
rect -1596 -143 -1592 -139
rect -1555 -143 -1551 -139
rect -1533 -143 -1529 -139
rect -1459 -143 -1455 -139
rect -1437 -143 -1433 -139
rect -1390 -143 -1386 -139
rect -380 -138 -376 -134
rect -251 -138 -247 -134
rect -1574 -199 -1570 -195
rect -445 -179 -441 -175
rect -437 -179 -433 -175
rect -396 -179 -392 -175
rect -1418 -199 -1414 -195
rect -1514 -208 -1510 -204
rect -1478 -208 -1474 -204
rect -364 -179 -360 -175
rect -348 -179 -344 -175
rect -321 -180 -317 -176
rect -267 -179 -263 -175
rect 16 -161 20 -157
rect 145 -161 149 -157
rect -235 -179 -231 -175
rect -219 -179 -215 -175
rect -192 -180 -188 -176
rect -56 -179 -52 -175
rect -48 -179 -44 -175
rect 0 -179 4 -175
rect -399 -229 -395 -225
rect -383 -212 -379 -208
rect -298 -235 -294 -231
rect -270 -212 -266 -208
rect -254 -212 -250 -208
rect -169 -235 -165 -231
rect -142 -235 -138 -231
rect -116 -209 -112 -205
rect 32 -179 36 -175
rect 48 -179 52 -175
rect 75 -180 79 -176
rect 129 -179 133 -175
rect 161 -179 165 -175
rect 177 -179 181 -175
rect 204 -180 208 -176
rect -35 -234 -31 -230
rect -3 -232 1 -228
rect 13 -212 17 -208
rect 98 -235 102 -231
rect -380 -281 -376 -277
rect -356 -281 -352 -277
rect -340 -281 -336 -277
rect -313 -280 -309 -276
rect 126 -212 130 -208
rect 142 -212 146 -208
rect 227 -235 231 -231
rect 254 -235 258 -231
rect 280 -209 284 -205
rect -251 -281 -247 -277
rect -227 -281 -223 -277
rect -211 -281 -207 -277
rect -184 -280 -180 -276
rect -131 -280 -127 -276
rect 16 -281 20 -277
rect 40 -281 44 -277
rect 56 -281 60 -277
rect 83 -280 87 -276
rect 145 -281 149 -277
rect 169 -281 173 -277
rect 185 -281 189 -277
rect 212 -280 216 -276
rect 265 -280 269 -276
rect -1574 -293 -1570 -289
rect -1418 -293 -1414 -289
rect -1514 -302 -1510 -298
rect -1478 -302 -1474 -298
rect -1615 -351 -1611 -347
rect -1596 -351 -1592 -347
rect -1555 -351 -1551 -347
rect -1533 -351 -1529 -347
rect -1459 -351 -1455 -347
rect -1437 -351 -1433 -347
rect -1390 -351 -1386 -347
rect -423 -344 -419 -340
rect -1574 -407 -1570 -403
rect -861 -386 -857 -382
rect -853 -386 -849 -382
rect -805 -386 -801 -382
rect -773 -386 -769 -382
rect -757 -386 -753 -382
rect -1418 -407 -1414 -403
rect -1514 -416 -1510 -412
rect -1478 -416 -1474 -412
rect -730 -387 -726 -383
rect -676 -386 -672 -382
rect -644 -386 -640 -382
rect -628 -386 -624 -382
rect -601 -387 -597 -383
rect -451 -386 -447 -382
rect -443 -386 -439 -382
rect -402 -386 -398 -382
rect -840 -441 -836 -437
rect -808 -439 -804 -435
rect -792 -419 -788 -415
rect -707 -442 -703 -438
rect -679 -419 -675 -415
rect -663 -419 -659 -415
rect -578 -442 -574 -438
rect -551 -442 -547 -438
rect -525 -416 -521 -412
rect -250 -346 -246 -342
rect -370 -386 -366 -382
rect -354 -386 -350 -382
rect -327 -387 -323 -383
rect -273 -386 -269 -382
rect 24 -364 28 -360
rect -241 -386 -237 -382
rect -225 -386 -221 -382
rect -198 -387 -194 -383
rect -405 -436 -401 -432
rect -389 -419 -385 -415
rect -304 -442 -300 -438
rect -789 -488 -785 -484
rect -765 -488 -761 -484
rect -749 -488 -745 -484
rect -722 -487 -718 -483
rect -276 -419 -272 -415
rect -260 -419 -256 -415
rect -175 -442 -171 -438
rect -148 -442 -144 -438
rect -122 -416 -118 -412
rect -660 -488 -656 -484
rect -636 -488 -632 -484
rect -620 -488 -616 -484
rect -593 -487 -589 -483
rect -540 -487 -536 -483
rect -386 -488 -382 -484
rect -362 -488 -358 -484
rect -346 -488 -342 -484
rect -319 -487 -315 -483
rect -257 -488 -253 -484
rect -233 -488 -229 -484
rect -217 -488 -213 -484
rect -190 -487 -186 -483
rect -137 -487 -133 -483
rect -1577 -516 -1573 -512
rect -1421 -516 -1417 -512
rect -1517 -525 -1513 -521
rect -1481 -525 -1477 -521
rect -1618 -574 -1614 -570
rect -1599 -574 -1595 -570
rect -1558 -574 -1554 -570
rect -1536 -574 -1532 -570
rect -1462 -574 -1458 -570
rect -1440 -574 -1436 -570
rect -1393 -574 -1389 -570
rect -1214 -566 -1210 -562
rect -1577 -630 -1573 -626
rect -1421 -630 -1417 -626
rect -1230 -630 -1226 -626
rect -1517 -639 -1513 -635
rect -1481 -639 -1477 -635
rect -1085 -604 -1081 -600
rect -1198 -630 -1194 -626
rect -1182 -630 -1178 -626
rect -1155 -631 -1151 -627
rect -1101 -630 -1097 -626
rect -1069 -630 -1065 -626
rect -1053 -630 -1049 -626
rect -1026 -631 -1022 -627
rect -850 -630 -846 -626
rect -293 -604 -289 -600
rect -818 -630 -814 -626
rect -802 -630 -798 -626
rect -775 -631 -771 -627
rect -721 -630 -717 -626
rect -689 -630 -685 -626
rect -673 -630 -669 -626
rect -646 -631 -642 -627
rect -1233 -663 -1229 -659
rect -1217 -663 -1213 -659
rect -1132 -686 -1128 -682
rect -1104 -663 -1100 -659
rect -1088 -663 -1084 -659
rect -1003 -686 -999 -682
rect -976 -686 -972 -682
rect -950 -660 -946 -656
rect -752 -686 -748 -682
rect -1214 -732 -1210 -728
rect -1190 -732 -1186 -728
rect -1174 -732 -1170 -728
rect -1147 -731 -1143 -727
rect -724 -663 -720 -659
rect -708 -663 -704 -659
rect -623 -686 -619 -682
rect -596 -686 -592 -682
rect -570 -660 -566 -656
rect -1085 -732 -1081 -728
rect -1061 -732 -1057 -728
rect -1045 -732 -1041 -728
rect -1018 -731 -1014 -727
rect -965 -731 -961 -727
rect -834 -732 -830 -728
rect -810 -732 -806 -728
rect -794 -732 -790 -728
rect -767 -731 -763 -727
rect -705 -732 -701 -728
rect -681 -732 -677 -728
rect -665 -732 -661 -728
rect -638 -731 -634 -727
rect -585 -731 -581 -727
rect -1177 -816 -1173 -812
rect -787 -813 -783 -809
rect -1158 -878 -1154 -874
rect -1002 -878 -998 -874
rect -1098 -887 -1094 -883
rect -1062 -887 -1058 -883
rect -768 -861 -764 -857
rect -612 -861 -608 -857
rect -708 -870 -704 -866
rect -672 -870 -668 -866
rect -276 -819 -272 -815
rect -276 -860 -272 -856
rect -120 -860 -116 -856
rect -216 -869 -212 -865
rect -180 -869 -176 -865
rect 116 -864 120 -860
rect -1199 -936 -1195 -932
rect -1139 -936 -1135 -932
rect -1117 -936 -1113 -932
rect -1043 -936 -1039 -932
rect -1021 -936 -1017 -932
rect -974 -936 -970 -932
rect -809 -919 -805 -915
rect -749 -919 -745 -915
rect -727 -919 -723 -915
rect -653 -919 -649 -915
rect -631 -919 -627 -915
rect -584 -919 -580 -915
rect -317 -918 -313 -914
rect -257 -918 -253 -914
rect -235 -918 -231 -914
rect -161 -918 -157 -914
rect -139 -918 -135 -914
rect -92 -918 -88 -914
rect 135 -875 139 -871
rect 291 -875 295 -871
rect 195 -884 199 -880
rect 231 -884 235 -880
rect 94 -933 98 -929
rect -1158 -992 -1154 -988
rect -768 -975 -764 -971
rect -612 -975 -608 -971
rect -276 -974 -272 -970
rect 154 -933 158 -929
rect 176 -933 180 -929
rect 250 -933 254 -929
rect 272 -933 276 -929
rect 319 -933 323 -929
rect -120 -974 -116 -970
rect -708 -984 -704 -980
rect -672 -984 -668 -980
rect -216 -983 -212 -979
rect -180 -983 -176 -979
rect -1002 -992 -998 -988
rect 135 -989 139 -985
rect 291 -989 295 -985
rect -1098 -1001 -1094 -997
rect -1062 -1001 -1058 -997
rect 195 -998 199 -994
rect 231 -998 235 -994
<< ndcontact >>
rect -1614 -6 -1610 -2
rect -1606 -6 -1602 -2
rect -1595 -6 -1591 -2
rect -1587 -6 -1583 -2
rect -1576 -6 -1572 -2
rect -1568 -6 -1564 -2
rect -1554 -6 -1550 2
rect -1546 -6 -1542 2
rect -1532 -6 -1528 -2
rect -1524 -6 -1520 -2
rect -1516 -6 -1512 -2
rect -1508 -6 -1504 -2
rect -1480 -6 -1476 -2
rect -1472 -6 -1468 -2
rect -1458 -6 -1454 2
rect -1450 -6 -1446 2
rect -1436 -6 -1432 -2
rect -1428 -6 -1424 -2
rect -1420 -6 -1416 -2
rect -1412 -6 -1408 -2
rect -1389 -6 -1385 -2
rect -1381 -6 -1377 -2
rect -1616 -162 -1612 -158
rect -1608 -162 -1604 -158
rect -1597 -162 -1593 -158
rect -1589 -162 -1585 -158
rect -1578 -162 -1574 -158
rect -1570 -162 -1566 -158
rect -1556 -162 -1552 -154
rect -1548 -162 -1544 -154
rect -1534 -162 -1530 -158
rect -1526 -162 -1522 -158
rect -1518 -162 -1514 -158
rect -1510 -162 -1506 -158
rect -1482 -162 -1478 -158
rect -1474 -162 -1470 -158
rect -1460 -162 -1456 -154
rect -1452 -162 -1448 -154
rect -1438 -162 -1434 -158
rect -1430 -162 -1426 -158
rect -1422 -162 -1418 -158
rect -1414 -162 -1410 -158
rect -1391 -162 -1387 -158
rect -1383 -162 -1379 -158
rect -449 -247 -445 -239
rect -433 -247 -429 -239
rect -400 -264 -396 -260
rect -392 -264 -388 -260
rect -384 -264 -380 -260
rect -376 -264 -372 -260
rect -368 -264 -364 -256
rect -352 -264 -348 -256
rect -336 -264 -332 -256
rect -327 -264 -323 -256
rect -307 -264 -303 -256
rect -299 -264 -295 -260
rect -291 -264 -287 -260
rect -271 -264 -267 -260
rect -263 -264 -259 -260
rect -255 -264 -251 -260
rect -247 -264 -243 -260
rect -239 -264 -235 -256
rect -223 -264 -219 -256
rect -207 -264 -203 -256
rect -198 -264 -194 -256
rect -178 -264 -174 -256
rect -170 -264 -166 -260
rect -162 -264 -158 -260
rect -144 -263 -140 -255
rect -135 -263 -131 -255
rect -127 -263 -123 -255
rect -60 -250 -56 -242
rect -44 -250 -40 -242
rect -36 -250 -32 -246
rect -28 -250 -24 -246
rect -118 -264 -114 -260
rect -108 -264 -104 -260
rect -4 -264 0 -260
rect 4 -264 8 -260
rect 12 -264 16 -260
rect 20 -264 24 -260
rect 28 -264 32 -256
rect 44 -264 48 -256
rect 60 -264 64 -256
rect 69 -264 73 -256
rect 89 -264 93 -256
rect 97 -264 101 -260
rect 105 -264 109 -260
rect 125 -264 129 -260
rect 133 -264 137 -260
rect 141 -264 145 -260
rect 149 -264 153 -260
rect 157 -264 161 -256
rect 173 -264 177 -256
rect 189 -264 193 -256
rect 198 -264 202 -256
rect 218 -264 222 -256
rect 226 -264 230 -260
rect 234 -264 238 -260
rect 252 -263 256 -255
rect 261 -263 265 -255
rect 269 -263 273 -255
rect 278 -264 282 -260
rect 288 -264 292 -260
rect -1616 -370 -1612 -366
rect -1608 -370 -1604 -366
rect -1597 -370 -1593 -366
rect -1589 -370 -1585 -366
rect -1578 -370 -1574 -366
rect -1570 -370 -1566 -366
rect -1556 -370 -1552 -362
rect -1548 -370 -1544 -362
rect -1534 -370 -1530 -366
rect -1526 -370 -1522 -366
rect -1518 -370 -1514 -366
rect -1510 -370 -1506 -366
rect -1482 -370 -1478 -366
rect -1474 -370 -1470 -366
rect -1460 -370 -1456 -362
rect -1452 -370 -1448 -362
rect -1438 -370 -1434 -366
rect -1430 -370 -1426 -366
rect -1422 -370 -1418 -366
rect -1414 -370 -1410 -366
rect -1391 -370 -1387 -366
rect -1383 -370 -1379 -366
rect -865 -457 -861 -449
rect -849 -457 -845 -449
rect -841 -457 -837 -453
rect -833 -457 -829 -453
rect -809 -471 -805 -467
rect -801 -471 -797 -467
rect -793 -471 -789 -467
rect -785 -471 -781 -467
rect -777 -471 -773 -463
rect -761 -471 -757 -463
rect -745 -471 -741 -463
rect -736 -471 -732 -463
rect -716 -471 -712 -463
rect -708 -471 -704 -467
rect -700 -471 -696 -467
rect -680 -471 -676 -467
rect -672 -471 -668 -467
rect -664 -471 -660 -467
rect -656 -471 -652 -467
rect -648 -471 -644 -463
rect -632 -471 -628 -463
rect -616 -471 -612 -463
rect -607 -471 -603 -463
rect -587 -471 -583 -463
rect -579 -471 -575 -467
rect -571 -471 -567 -467
rect -553 -470 -549 -462
rect -544 -470 -540 -462
rect -536 -470 -532 -462
rect -455 -454 -451 -446
rect -439 -454 -435 -446
rect -527 -471 -523 -467
rect -517 -471 -513 -467
rect -406 -471 -402 -467
rect -398 -471 -394 -467
rect -390 -471 -386 -467
rect -382 -471 -378 -467
rect -374 -471 -370 -463
rect -358 -471 -354 -463
rect -342 -471 -338 -463
rect -333 -471 -329 -463
rect -313 -471 -309 -463
rect -305 -471 -301 -467
rect -297 -471 -293 -467
rect -277 -471 -273 -467
rect -269 -471 -265 -467
rect -261 -471 -257 -467
rect -253 -471 -249 -467
rect -245 -471 -241 -463
rect -229 -471 -225 -463
rect -213 -471 -209 -463
rect -204 -471 -200 -463
rect -184 -471 -180 -463
rect -176 -471 -172 -467
rect -168 -471 -164 -467
rect -150 -470 -146 -462
rect -141 -470 -137 -462
rect -133 -470 -129 -462
rect -124 -471 -120 -467
rect -114 -471 -110 -467
rect -1619 -593 -1615 -589
rect -1611 -593 -1607 -589
rect -1600 -593 -1596 -589
rect -1592 -593 -1588 -589
rect -1581 -593 -1577 -589
rect -1573 -593 -1569 -589
rect -1559 -593 -1555 -585
rect -1551 -593 -1547 -585
rect -1537 -593 -1533 -589
rect -1529 -593 -1525 -589
rect -1521 -593 -1517 -589
rect -1513 -593 -1509 -589
rect -1485 -593 -1481 -589
rect -1477 -593 -1473 -589
rect -1463 -593 -1459 -585
rect -1455 -593 -1451 -585
rect -1441 -593 -1437 -589
rect -1433 -593 -1429 -589
rect -1425 -593 -1421 -589
rect -1417 -593 -1413 -589
rect -1394 -593 -1390 -589
rect -1386 -593 -1382 -589
rect -1234 -715 -1230 -711
rect -1226 -715 -1222 -711
rect -1218 -715 -1214 -711
rect -1210 -715 -1206 -711
rect -1202 -715 -1198 -707
rect -1186 -715 -1182 -707
rect -1170 -715 -1166 -707
rect -1161 -715 -1157 -707
rect -1141 -715 -1137 -707
rect -1133 -715 -1129 -711
rect -1125 -715 -1121 -711
rect -1105 -715 -1101 -711
rect -1097 -715 -1093 -711
rect -1089 -715 -1085 -711
rect -1081 -715 -1077 -711
rect -1073 -715 -1069 -707
rect -1057 -715 -1053 -707
rect -1041 -715 -1037 -707
rect -1032 -715 -1028 -707
rect -1012 -715 -1008 -707
rect -1004 -715 -1000 -711
rect -996 -715 -992 -711
rect -978 -714 -974 -706
rect -969 -714 -965 -706
rect -961 -714 -957 -706
rect -952 -715 -948 -711
rect -942 -715 -938 -711
rect -854 -715 -850 -711
rect -846 -715 -842 -711
rect -838 -715 -834 -711
rect -830 -715 -826 -711
rect -822 -715 -818 -707
rect -806 -715 -802 -707
rect -790 -715 -786 -707
rect -781 -715 -777 -707
rect -761 -715 -757 -707
rect -753 -715 -749 -711
rect -745 -715 -741 -711
rect -725 -715 -721 -711
rect -717 -715 -713 -711
rect -709 -715 -705 -711
rect -701 -715 -697 -711
rect -693 -715 -689 -707
rect -677 -715 -673 -707
rect -661 -715 -657 -707
rect -652 -715 -648 -707
rect -632 -715 -628 -707
rect -624 -715 -620 -711
rect -616 -715 -612 -711
rect -598 -714 -594 -706
rect -589 -714 -585 -706
rect -581 -714 -577 -706
rect -572 -715 -568 -711
rect -562 -715 -558 -711
rect -1200 -955 -1196 -951
rect -1192 -955 -1188 -951
rect -1181 -955 -1177 -951
rect -1173 -955 -1169 -951
rect -1162 -955 -1158 -951
rect -1154 -955 -1150 -951
rect -1140 -955 -1136 -947
rect -1132 -955 -1128 -947
rect -1118 -955 -1114 -951
rect -1110 -955 -1106 -951
rect -1102 -955 -1098 -951
rect -1094 -955 -1090 -951
rect -1066 -955 -1062 -951
rect -1058 -955 -1054 -951
rect -1044 -955 -1040 -947
rect -1036 -955 -1032 -947
rect -810 -938 -806 -934
rect -802 -938 -798 -934
rect -791 -938 -787 -934
rect -783 -938 -779 -934
rect -772 -938 -768 -934
rect -764 -938 -760 -934
rect -750 -938 -746 -930
rect -742 -938 -738 -930
rect -728 -938 -724 -934
rect -720 -938 -716 -934
rect -712 -938 -708 -934
rect -704 -938 -700 -934
rect -676 -938 -672 -934
rect -668 -938 -664 -934
rect -654 -938 -650 -930
rect -646 -938 -642 -930
rect -632 -938 -628 -934
rect -624 -938 -620 -934
rect -616 -938 -612 -934
rect -608 -938 -604 -934
rect -585 -938 -581 -934
rect -577 -938 -573 -934
rect -318 -937 -314 -933
rect -310 -937 -306 -933
rect -299 -937 -295 -933
rect -291 -937 -287 -933
rect -280 -937 -276 -933
rect -272 -937 -268 -933
rect -258 -937 -254 -929
rect -250 -937 -246 -929
rect -236 -937 -232 -933
rect -228 -937 -224 -933
rect -220 -937 -216 -933
rect -212 -937 -208 -933
rect -184 -937 -180 -933
rect -176 -937 -172 -933
rect -162 -937 -158 -929
rect -154 -937 -150 -929
rect -140 -937 -136 -933
rect -132 -937 -128 -933
rect -124 -937 -120 -933
rect -116 -937 -112 -933
rect -93 -937 -89 -933
rect -85 -937 -81 -933
rect -1022 -955 -1018 -951
rect -1014 -955 -1010 -951
rect -1006 -955 -1002 -951
rect -998 -955 -994 -951
rect -975 -955 -971 -951
rect -967 -955 -963 -951
rect 93 -952 97 -948
rect 101 -952 105 -948
rect 112 -952 116 -948
rect 120 -952 124 -948
rect 131 -952 135 -948
rect 139 -952 143 -948
rect 153 -952 157 -944
rect 161 -952 165 -944
rect 175 -952 179 -948
rect 183 -952 187 -948
rect 191 -952 195 -948
rect 199 -952 203 -948
rect 227 -952 231 -948
rect 235 -952 239 -948
rect 249 -952 253 -944
rect 257 -952 261 -944
rect 271 -952 275 -948
rect 279 -952 283 -948
rect 287 -952 291 -948
rect 295 -952 299 -948
rect 318 -952 322 -948
rect 326 -952 330 -948
<< pdcontact >>
rect -1614 33 -1610 41
rect -1606 33 -1602 41
rect -1595 33 -1591 41
rect -1587 33 -1583 41
rect -1576 33 -1572 41
rect -1568 33 -1564 41
rect -1554 25 -1550 41
rect -1546 25 -1542 41
rect -1532 33 -1528 41
rect -1524 33 -1520 41
rect -1516 33 -1512 41
rect -1508 33 -1504 41
rect -1480 33 -1476 41
rect -1472 33 -1468 41
rect -1458 25 -1454 41
rect -1450 25 -1446 41
rect -1436 33 -1432 41
rect -1428 33 -1424 41
rect -1420 33 -1416 41
rect -1412 33 -1408 41
rect -1389 33 -1385 41
rect -1381 33 -1377 41
rect -1616 -123 -1612 -115
rect -1608 -123 -1604 -115
rect -1597 -123 -1593 -115
rect -1589 -123 -1585 -115
rect -1578 -123 -1574 -115
rect -1570 -123 -1566 -115
rect -1556 -131 -1552 -115
rect -1548 -131 -1544 -115
rect -1534 -123 -1530 -115
rect -1526 -123 -1522 -115
rect -1518 -123 -1514 -115
rect -1510 -123 -1506 -115
rect -1482 -123 -1478 -115
rect -1474 -123 -1470 -115
rect -1460 -131 -1456 -115
rect -1452 -131 -1448 -115
rect -1438 -123 -1434 -115
rect -1430 -123 -1426 -115
rect -1422 -123 -1418 -115
rect -1414 -123 -1410 -115
rect -1391 -123 -1387 -115
rect -1383 -123 -1379 -115
rect -400 -200 -396 -192
rect -392 -200 -388 -192
rect -384 -200 -380 -192
rect -376 -200 -372 -192
rect -449 -213 -445 -205
rect -441 -213 -437 -205
rect -433 -213 -429 -205
rect -368 -208 -364 -192
rect -360 -200 -356 -192
rect -352 -208 -348 -192
rect -344 -208 -340 -200
rect -336 -208 -332 -192
rect -326 -198 -322 -194
rect -317 -198 -313 -194
rect -308 -198 -304 -194
rect -299 -200 -295 -192
rect -291 -200 -287 -192
rect -271 -200 -267 -192
rect -263 -200 -259 -192
rect -255 -200 -251 -192
rect -247 -200 -243 -192
rect -239 -208 -235 -192
rect -231 -200 -227 -192
rect -223 -208 -219 -192
rect -215 -208 -211 -200
rect -207 -208 -203 -192
rect -197 -198 -193 -194
rect -188 -198 -184 -194
rect -179 -198 -175 -194
rect -170 -200 -166 -192
rect -162 -200 -158 -192
rect -144 -200 -140 -192
rect -127 -200 -123 -192
rect -118 -200 -114 -192
rect -108 -200 -104 -192
rect -4 -200 0 -192
rect 4 -200 8 -192
rect 12 -200 16 -192
rect 20 -200 24 -192
rect -60 -216 -56 -208
rect -52 -216 -48 -208
rect -44 -216 -40 -208
rect -36 -216 -32 -208
rect -28 -216 -24 -208
rect 28 -208 32 -192
rect 36 -200 40 -192
rect 44 -208 48 -192
rect 52 -208 56 -200
rect 60 -208 64 -192
rect 70 -198 74 -194
rect 79 -198 83 -194
rect 88 -198 92 -194
rect 97 -200 101 -192
rect 105 -200 109 -192
rect 125 -200 129 -192
rect 133 -200 137 -192
rect 141 -200 145 -192
rect 149 -200 153 -192
rect 157 -208 161 -192
rect 165 -200 169 -192
rect 173 -208 177 -192
rect 181 -208 185 -200
rect 189 -208 193 -192
rect 199 -198 203 -194
rect 208 -198 212 -194
rect 217 -198 221 -194
rect 226 -200 230 -192
rect 234 -200 238 -192
rect 252 -200 256 -192
rect 269 -200 273 -192
rect 278 -200 282 -192
rect 288 -200 292 -192
rect -1616 -331 -1612 -323
rect -1608 -331 -1604 -323
rect -1597 -331 -1593 -323
rect -1589 -331 -1585 -323
rect -1578 -331 -1574 -323
rect -1570 -331 -1566 -323
rect -1556 -339 -1552 -323
rect -1548 -339 -1544 -323
rect -1534 -331 -1530 -323
rect -1526 -331 -1522 -323
rect -1518 -331 -1514 -323
rect -1510 -331 -1506 -323
rect -1482 -331 -1478 -323
rect -1474 -331 -1470 -323
rect -1460 -339 -1456 -323
rect -1452 -339 -1448 -323
rect -1438 -331 -1434 -323
rect -1430 -331 -1426 -323
rect -1422 -331 -1418 -323
rect -1414 -331 -1410 -323
rect -1391 -331 -1387 -323
rect -1383 -331 -1379 -323
rect -809 -407 -805 -399
rect -801 -407 -797 -399
rect -793 -407 -789 -399
rect -785 -407 -781 -399
rect -865 -423 -861 -415
rect -857 -423 -853 -415
rect -849 -423 -845 -415
rect -841 -423 -837 -415
rect -833 -423 -829 -415
rect -777 -415 -773 -399
rect -769 -407 -765 -399
rect -761 -415 -757 -399
rect -753 -415 -749 -407
rect -745 -415 -741 -399
rect -735 -405 -731 -401
rect -726 -405 -722 -401
rect -717 -405 -713 -401
rect -708 -407 -704 -399
rect -700 -407 -696 -399
rect -680 -407 -676 -399
rect -672 -407 -668 -399
rect -664 -407 -660 -399
rect -656 -407 -652 -399
rect -648 -415 -644 -399
rect -640 -407 -636 -399
rect -632 -415 -628 -399
rect -624 -415 -620 -407
rect -616 -415 -612 -399
rect -606 -405 -602 -401
rect -597 -405 -593 -401
rect -588 -405 -584 -401
rect -579 -407 -575 -399
rect -571 -407 -567 -399
rect -553 -407 -549 -399
rect -536 -407 -532 -399
rect -527 -407 -523 -399
rect -517 -407 -513 -399
rect -406 -407 -402 -399
rect -398 -407 -394 -399
rect -390 -407 -386 -399
rect -382 -407 -378 -399
rect -455 -420 -451 -412
rect -447 -420 -443 -412
rect -439 -420 -435 -412
rect -374 -415 -370 -399
rect -366 -407 -362 -399
rect -358 -415 -354 -399
rect -350 -415 -346 -407
rect -342 -415 -338 -399
rect -332 -405 -328 -401
rect -323 -405 -319 -401
rect -314 -405 -310 -401
rect -305 -407 -301 -399
rect -297 -407 -293 -399
rect -277 -407 -273 -399
rect -269 -407 -265 -399
rect -261 -407 -257 -399
rect -253 -407 -249 -399
rect -245 -415 -241 -399
rect -237 -407 -233 -399
rect -229 -415 -225 -399
rect -221 -415 -217 -407
rect -213 -415 -209 -399
rect -203 -405 -199 -401
rect -194 -405 -190 -401
rect -185 -405 -181 -401
rect -176 -407 -172 -399
rect -168 -407 -164 -399
rect -150 -407 -146 -399
rect -133 -407 -129 -399
rect -124 -407 -120 -399
rect -114 -407 -110 -399
rect -1619 -554 -1615 -546
rect -1611 -554 -1607 -546
rect -1600 -554 -1596 -546
rect -1592 -554 -1588 -546
rect -1581 -554 -1577 -546
rect -1573 -554 -1569 -546
rect -1559 -562 -1555 -546
rect -1551 -562 -1547 -546
rect -1537 -554 -1533 -546
rect -1529 -554 -1525 -546
rect -1521 -554 -1517 -546
rect -1513 -554 -1509 -546
rect -1485 -554 -1481 -546
rect -1477 -554 -1473 -546
rect -1463 -562 -1459 -546
rect -1455 -562 -1451 -546
rect -1441 -554 -1437 -546
rect -1433 -554 -1429 -546
rect -1425 -554 -1421 -546
rect -1417 -554 -1413 -546
rect -1394 -554 -1390 -546
rect -1386 -554 -1382 -546
rect -1234 -651 -1230 -643
rect -1226 -651 -1222 -643
rect -1218 -651 -1214 -643
rect -1210 -651 -1206 -643
rect -1202 -659 -1198 -643
rect -1194 -651 -1190 -643
rect -1186 -659 -1182 -643
rect -1178 -659 -1174 -651
rect -1170 -659 -1166 -643
rect -1160 -649 -1156 -645
rect -1151 -649 -1147 -645
rect -1142 -649 -1138 -645
rect -1133 -651 -1129 -643
rect -1125 -651 -1121 -643
rect -1105 -651 -1101 -643
rect -1097 -651 -1093 -643
rect -1089 -651 -1085 -643
rect -1081 -651 -1077 -643
rect -1073 -659 -1069 -643
rect -1065 -651 -1061 -643
rect -1057 -659 -1053 -643
rect -1049 -659 -1045 -651
rect -1041 -659 -1037 -643
rect -1031 -649 -1027 -645
rect -1022 -649 -1018 -645
rect -1013 -649 -1009 -645
rect -1004 -651 -1000 -643
rect -996 -651 -992 -643
rect -978 -651 -974 -643
rect -961 -651 -957 -643
rect -952 -651 -948 -643
rect -942 -651 -938 -643
rect -854 -651 -850 -643
rect -846 -651 -842 -643
rect -838 -651 -834 -643
rect -830 -651 -826 -643
rect -822 -659 -818 -643
rect -814 -651 -810 -643
rect -806 -659 -802 -643
rect -798 -659 -794 -651
rect -790 -659 -786 -643
rect -780 -649 -776 -645
rect -771 -649 -767 -645
rect -762 -649 -758 -645
rect -753 -651 -749 -643
rect -745 -651 -741 -643
rect -725 -651 -721 -643
rect -717 -651 -713 -643
rect -709 -651 -705 -643
rect -701 -651 -697 -643
rect -693 -659 -689 -643
rect -685 -651 -681 -643
rect -677 -659 -673 -643
rect -669 -659 -665 -651
rect -661 -659 -657 -643
rect -651 -649 -647 -645
rect -642 -649 -638 -645
rect -633 -649 -629 -645
rect -624 -651 -620 -643
rect -616 -651 -612 -643
rect -598 -651 -594 -643
rect -581 -651 -577 -643
rect -572 -651 -568 -643
rect -562 -651 -558 -643
rect -810 -899 -806 -891
rect -802 -899 -798 -891
rect -791 -899 -787 -891
rect -783 -899 -779 -891
rect -772 -899 -768 -891
rect -764 -899 -760 -891
rect -1200 -916 -1196 -908
rect -1192 -916 -1188 -908
rect -1181 -916 -1177 -908
rect -1173 -916 -1169 -908
rect -1162 -916 -1158 -908
rect -1154 -916 -1150 -908
rect -1140 -924 -1136 -908
rect -1132 -924 -1128 -908
rect -1118 -916 -1114 -908
rect -1110 -916 -1106 -908
rect -1102 -916 -1098 -908
rect -1094 -916 -1090 -908
rect -1066 -916 -1062 -908
rect -1058 -916 -1054 -908
rect -1044 -924 -1040 -908
rect -1036 -924 -1032 -908
rect -1022 -916 -1018 -908
rect -1014 -916 -1010 -908
rect -1006 -916 -1002 -908
rect -998 -916 -994 -908
rect -975 -916 -971 -908
rect -967 -916 -963 -908
rect -750 -907 -746 -891
rect -742 -907 -738 -891
rect -728 -899 -724 -891
rect -720 -899 -716 -891
rect -712 -899 -708 -891
rect -704 -899 -700 -891
rect -676 -899 -672 -891
rect -668 -899 -664 -891
rect -654 -907 -650 -891
rect -646 -907 -642 -891
rect -632 -899 -628 -891
rect -624 -899 -620 -891
rect -616 -899 -612 -891
rect -608 -899 -604 -891
rect -585 -899 -581 -891
rect -577 -899 -573 -891
rect -318 -898 -314 -890
rect -310 -898 -306 -890
rect -299 -898 -295 -890
rect -291 -898 -287 -890
rect -280 -898 -276 -890
rect -272 -898 -268 -890
rect -258 -906 -254 -890
rect -250 -906 -246 -890
rect -236 -898 -232 -890
rect -228 -898 -224 -890
rect -220 -898 -216 -890
rect -212 -898 -208 -890
rect -184 -898 -180 -890
rect -176 -898 -172 -890
rect -162 -906 -158 -890
rect -154 -906 -150 -890
rect -140 -898 -136 -890
rect -132 -898 -128 -890
rect -124 -898 -120 -890
rect -116 -898 -112 -890
rect -93 -898 -89 -890
rect -85 -898 -81 -890
rect 93 -913 97 -905
rect 101 -913 105 -905
rect 112 -913 116 -905
rect 120 -913 124 -905
rect 131 -913 135 -905
rect 139 -913 143 -905
rect 153 -921 157 -905
rect 161 -921 165 -905
rect 175 -913 179 -905
rect 183 -913 187 -905
rect 191 -913 195 -905
rect 199 -913 203 -905
rect 227 -913 231 -905
rect 235 -913 239 -905
rect 249 -921 253 -905
rect 257 -921 261 -905
rect 271 -913 275 -905
rect 279 -913 283 -905
rect 287 -913 291 -905
rect 295 -913 299 -905
rect 318 -913 322 -905
rect 326 -913 330 -905
<< m2contact >>
rect -1605 61 -1600 66
rect -1606 13 -1601 18
rect -1568 13 -1563 18
rect -1539 13 -1535 17
rect -1508 13 -1503 18
rect -1481 13 -1476 18
rect -1464 13 -1459 18
rect -1443 13 -1438 18
rect -1412 13 -1407 18
rect -1398 13 -1393 18
rect -1373 13 -1369 17
rect -1605 -43 -1600 -38
rect -1624 -56 -1620 -52
rect -1624 -81 -1620 -77
rect -1607 -95 -1602 -90
rect -517 9 -513 13
rect -1608 -143 -1603 -138
rect -1570 -143 -1565 -138
rect -1541 -143 -1537 -139
rect -1510 -143 -1505 -138
rect -1483 -143 -1478 -138
rect -1466 -143 -1461 -138
rect -1445 -143 -1440 -138
rect -1414 -143 -1409 -138
rect -1400 -143 -1395 -138
rect -1375 -143 -1371 -139
rect -1607 -199 -1602 -194
rect -1626 -212 -1622 -208
rect -1626 -289 -1622 -285
rect -1607 -303 -1602 -298
rect -1608 -351 -1603 -346
rect -1570 -351 -1565 -346
rect -1541 -351 -1537 -347
rect -1510 -351 -1505 -346
rect -1483 -351 -1478 -346
rect -1466 -351 -1461 -346
rect -1445 -351 -1440 -346
rect -1414 -351 -1409 -346
rect -1400 -351 -1395 -346
rect -1375 -351 -1371 -347
rect -1607 -407 -1602 -402
rect -1626 -420 -1622 -416
rect -853 -147 -849 -143
rect -861 -379 -857 -375
rect -445 -156 -441 -152
rect -437 -172 -433 -168
rect -356 -179 -351 -174
rect -227 -179 -222 -174
rect 153 -161 157 -157
rect -48 -172 -44 -168
rect 40 -179 45 -174
rect 169 -179 174 -174
rect -392 -233 -387 -228
rect -376 -233 -371 -228
rect -332 -227 -327 -222
rect -277 -213 -272 -208
rect -284 -236 -279 -231
rect -263 -233 -258 -228
rect -247 -233 -242 -228
rect -203 -227 -198 -222
rect -77 -213 -73 -209
rect 4 -233 9 -228
rect 20 -233 25 -228
rect 64 -227 69 -222
rect 119 -213 124 -208
rect 112 -236 117 -231
rect 133 -233 138 -228
rect 149 -233 154 -228
rect 193 -227 198 -222
rect 295 -267 299 -263
rect -348 -282 -343 -277
rect -219 -282 -214 -277
rect -132 -287 -127 -282
rect 48 -282 53 -277
rect -103 -294 -99 -290
rect 177 -282 182 -277
rect 264 -287 269 -282
rect 336 -280 340 -276
rect -765 -386 -760 -381
rect -636 -386 -631 -381
rect -451 -379 -447 -375
rect -423 -338 -419 -334
rect 32 -364 36 -360
rect -362 -386 -357 -381
rect -233 -386 -228 -381
rect -1626 -512 -1622 -508
rect -1610 -526 -1605 -521
rect -801 -440 -796 -435
rect -785 -440 -780 -435
rect -741 -434 -736 -429
rect -686 -420 -681 -415
rect -693 -443 -688 -438
rect -672 -440 -667 -435
rect -656 -440 -651 -435
rect -612 -434 -607 -429
rect -508 -455 -504 -451
rect -398 -440 -393 -435
rect -382 -440 -377 -435
rect -338 -434 -333 -429
rect -283 -420 -278 -415
rect -290 -443 -285 -438
rect -269 -440 -264 -435
rect -253 -440 -248 -435
rect -209 -434 -204 -429
rect -106 -468 -102 -464
rect -757 -489 -752 -484
rect -628 -489 -623 -484
rect -541 -494 -536 -489
rect -354 -489 -349 -484
rect -225 -489 -220 -484
rect -138 -494 -133 -489
rect -1611 -574 -1606 -569
rect -1573 -574 -1568 -569
rect -1544 -574 -1540 -570
rect -1513 -574 -1508 -569
rect -1486 -574 -1481 -569
rect -1469 -574 -1464 -569
rect -1448 -574 -1443 -569
rect -1417 -574 -1412 -569
rect -1403 -574 -1398 -569
rect -1378 -574 -1374 -570
rect -1610 -630 -1605 -625
rect -1626 -643 -1622 -639
rect -1214 -558 -1210 -554
rect -1190 -630 -1185 -625
rect -1061 -630 -1056 -625
rect -850 -622 -846 -618
rect -810 -630 -805 -625
rect -681 -630 -676 -625
rect -1226 -684 -1221 -679
rect -1210 -684 -1205 -679
rect -1166 -678 -1161 -673
rect -1111 -664 -1106 -659
rect -1118 -687 -1113 -682
rect -1097 -684 -1092 -679
rect -1081 -684 -1076 -679
rect -1037 -678 -1032 -673
rect -846 -684 -841 -679
rect -830 -684 -825 -679
rect -786 -678 -781 -673
rect -731 -664 -726 -659
rect -738 -687 -733 -682
rect -717 -684 -712 -679
rect -701 -684 -696 -679
rect -657 -678 -652 -673
rect -285 -604 -281 -600
rect -1182 -733 -1177 -728
rect -1053 -733 -1048 -728
rect -966 -738 -961 -733
rect -802 -733 -797 -728
rect -673 -733 -668 -728
rect -586 -738 -581 -733
rect -1169 -816 -1165 -812
rect -780 -813 -776 -809
rect -268 -819 -264 -815
rect -1191 -888 -1186 -883
rect -1192 -936 -1187 -931
rect -1154 -936 -1149 -931
rect -1125 -936 -1121 -932
rect -1094 -936 -1089 -931
rect -1067 -936 -1062 -931
rect -1050 -936 -1045 -931
rect -1029 -936 -1024 -931
rect -998 -936 -993 -931
rect -984 -936 -979 -931
rect -801 -871 -796 -866
rect -802 -919 -797 -914
rect -1191 -992 -1186 -987
rect -1210 -1006 -1206 -1001
rect -764 -919 -759 -914
rect -735 -919 -731 -915
rect -704 -919 -699 -914
rect -677 -919 -672 -914
rect -660 -919 -655 -914
rect -639 -919 -634 -914
rect -608 -919 -603 -914
rect -594 -919 -589 -914
rect -309 -870 -304 -865
rect 124 -864 128 -860
rect -310 -918 -305 -913
rect -801 -975 -796 -970
rect -811 -988 -807 -984
rect -272 -918 -267 -913
rect -243 -918 -239 -914
rect -212 -918 -207 -913
rect -185 -918 -180 -913
rect -168 -918 -163 -913
rect -147 -918 -142 -913
rect -116 -918 -111 -913
rect -102 -918 -97 -913
rect 102 -885 107 -880
rect 101 -933 106 -928
rect -309 -974 -304 -969
rect -323 -987 -319 -983
rect 139 -933 144 -928
rect 168 -933 172 -929
rect 199 -933 204 -928
rect 226 -933 231 -928
rect 243 -933 248 -928
rect 264 -933 269 -928
rect 295 -933 300 -928
rect 309 -933 314 -928
rect 102 -989 107 -984
rect 87 -1002 91 -998
<< psubstratepcontact >>
rect -1613 -14 -1609 -10
rect -1594 -14 -1590 -10
rect -1553 -14 -1549 -10
rect -1531 -14 -1527 -10
rect -1457 -14 -1453 -10
rect -1435 -14 -1431 -10
rect -1388 -14 -1384 -10
rect -1615 -170 -1611 -166
rect -1596 -170 -1592 -166
rect -1555 -170 -1551 -166
rect -1533 -170 -1529 -166
rect -1459 -170 -1455 -166
rect -1437 -170 -1433 -166
rect -1390 -170 -1386 -166
rect -448 -272 -444 -268
rect -399 -272 -395 -268
rect -326 -272 -322 -268
rect -308 -272 -304 -268
rect -298 -272 -294 -268
rect -270 -272 -266 -268
rect -197 -272 -193 -268
rect -179 -272 -175 -268
rect -169 -272 -165 -268
rect -136 -272 -132 -268
rect -118 -272 -114 -268
rect -59 -272 -55 -268
rect -35 -272 -31 -268
rect -3 -272 1 -268
rect 70 -272 74 -268
rect 88 -272 92 -268
rect 98 -272 102 -268
rect 126 -272 130 -268
rect 199 -272 203 -268
rect 217 -272 221 -268
rect 227 -272 231 -268
rect 260 -272 264 -268
rect 278 -272 282 -268
rect -1615 -378 -1611 -374
rect -1596 -378 -1592 -374
rect -1555 -378 -1551 -374
rect -1533 -378 -1529 -374
rect -1459 -378 -1455 -374
rect -1437 -378 -1433 -374
rect -1390 -378 -1386 -374
rect -864 -479 -860 -475
rect -840 -479 -836 -475
rect -808 -479 -804 -475
rect -735 -479 -731 -475
rect -717 -479 -713 -475
rect -707 -479 -703 -475
rect -679 -479 -675 -475
rect -606 -479 -602 -475
rect -588 -479 -584 -475
rect -578 -479 -574 -475
rect -545 -479 -541 -475
rect -527 -479 -523 -475
rect -454 -479 -450 -475
rect -405 -479 -401 -475
rect -332 -479 -328 -475
rect -314 -479 -310 -475
rect -304 -479 -300 -475
rect -276 -479 -272 -475
rect -203 -479 -199 -475
rect -185 -479 -181 -475
rect -175 -479 -171 -475
rect -142 -479 -138 -475
rect -124 -479 -120 -475
rect -1618 -601 -1614 -597
rect -1599 -601 -1595 -597
rect -1558 -601 -1554 -597
rect -1536 -601 -1532 -597
rect -1462 -601 -1458 -597
rect -1440 -601 -1436 -597
rect -1393 -601 -1389 -597
rect -1233 -723 -1229 -719
rect -1160 -723 -1156 -719
rect -1142 -723 -1138 -719
rect -1132 -723 -1128 -719
rect -1104 -723 -1100 -719
rect -1031 -723 -1027 -719
rect -1013 -723 -1009 -719
rect -1003 -723 -999 -719
rect -970 -723 -966 -719
rect -952 -723 -948 -719
rect -853 -723 -849 -719
rect -780 -723 -776 -719
rect -762 -723 -758 -719
rect -752 -723 -748 -719
rect -724 -723 -720 -719
rect -651 -723 -647 -719
rect -633 -723 -629 -719
rect -623 -723 -619 -719
rect -590 -723 -586 -719
rect -572 -723 -568 -719
rect -809 -946 -805 -942
rect -790 -946 -786 -942
rect -1199 -963 -1195 -959
rect -1180 -963 -1176 -959
rect -1139 -963 -1135 -959
rect -1117 -963 -1113 -959
rect -1043 -963 -1039 -959
rect -1021 -963 -1017 -959
rect -974 -963 -970 -959
rect -749 -946 -745 -942
rect -727 -946 -723 -942
rect -653 -946 -649 -942
rect -631 -946 -627 -942
rect -584 -946 -580 -942
rect -317 -945 -313 -941
rect -298 -945 -294 -941
rect -257 -945 -253 -941
rect -235 -945 -231 -941
rect -161 -945 -157 -941
rect -139 -945 -135 -941
rect -92 -945 -88 -941
rect 94 -960 98 -956
rect 113 -960 117 -956
rect 154 -960 158 -956
rect 176 -960 180 -956
rect 250 -960 254 -956
rect 272 -960 276 -956
rect 319 -960 323 -956
<< nsubstratencontact >>
rect -1613 45 -1609 49
rect -1594 45 -1590 49
rect -1553 45 -1549 49
rect -1531 45 -1527 49
rect -1457 45 -1453 49
rect -1435 45 -1431 49
rect -1388 45 -1384 49
rect -1615 -111 -1611 -107
rect -1596 -111 -1592 -107
rect -1555 -111 -1551 -107
rect -1533 -111 -1529 -107
rect -1459 -111 -1455 -107
rect -1437 -111 -1433 -107
rect -1390 -111 -1386 -107
rect -441 -188 -437 -184
rect -384 -188 -380 -184
rect -325 -188 -321 -184
rect -308 -188 -304 -184
rect -255 -188 -251 -184
rect -196 -188 -192 -184
rect -179 -188 -175 -184
rect -143 -188 -139 -184
rect -118 -188 -114 -184
rect -52 -188 -48 -184
rect -35 -188 -31 -184
rect 12 -188 16 -184
rect 71 -188 75 -184
rect 88 -188 92 -184
rect 141 -188 145 -184
rect 200 -188 204 -184
rect 217 -188 221 -184
rect 253 -188 257 -184
rect 278 -188 282 -184
rect -1615 -319 -1611 -315
rect -1596 -319 -1592 -315
rect -1555 -319 -1551 -315
rect -1533 -319 -1529 -315
rect -1459 -319 -1455 -315
rect -1437 -319 -1433 -315
rect -1390 -319 -1386 -315
rect -857 -395 -853 -391
rect -840 -395 -836 -391
rect -792 -395 -788 -391
rect -734 -395 -730 -391
rect -717 -395 -713 -391
rect -664 -395 -660 -391
rect -605 -395 -601 -391
rect -588 -395 -584 -391
rect -552 -395 -548 -391
rect -527 -395 -523 -391
rect -447 -395 -443 -391
rect -390 -395 -386 -391
rect -331 -395 -327 -391
rect -314 -395 -310 -391
rect -261 -395 -257 -391
rect -202 -395 -198 -391
rect -185 -395 -181 -391
rect -149 -395 -145 -391
rect -124 -395 -120 -391
rect -1618 -542 -1614 -538
rect -1599 -542 -1595 -538
rect -1558 -542 -1554 -538
rect -1536 -542 -1532 -538
rect -1462 -542 -1458 -538
rect -1440 -542 -1436 -538
rect -1393 -542 -1389 -538
rect -1218 -639 -1214 -635
rect -1159 -639 -1155 -635
rect -1142 -639 -1138 -635
rect -1089 -639 -1085 -635
rect -1030 -639 -1026 -635
rect -1013 -639 -1009 -635
rect -977 -639 -973 -635
rect -952 -639 -948 -635
rect -838 -639 -834 -635
rect -779 -639 -775 -635
rect -762 -639 -758 -635
rect -709 -639 -705 -635
rect -650 -639 -646 -635
rect -633 -639 -629 -635
rect -597 -639 -593 -635
rect -572 -639 -568 -635
rect -1199 -904 -1195 -900
rect -1181 -904 -1177 -900
rect -1139 -904 -1135 -900
rect -1117 -904 -1113 -900
rect -1043 -904 -1039 -900
rect -1021 -904 -1017 -900
rect -809 -887 -805 -883
rect -791 -887 -787 -883
rect -749 -887 -745 -883
rect -727 -887 -723 -883
rect -653 -887 -649 -883
rect -631 -887 -627 -883
rect -584 -887 -580 -883
rect -317 -886 -313 -882
rect -299 -886 -295 -882
rect -257 -886 -253 -882
rect -235 -886 -231 -882
rect -161 -886 -157 -882
rect -139 -886 -135 -882
rect -92 -886 -88 -882
rect -974 -904 -970 -900
rect 94 -901 98 -897
rect 112 -901 116 -897
rect 154 -901 158 -897
rect 176 -901 180 -897
rect 250 -901 254 -897
rect 272 -901 276 -897
rect 319 -901 323 -897
<< labels >>
rlabel metal1 -852 115 -852 115 1 vdd
rlabel metal1 -1731 -387 -1731 -387 3 gnd
rlabel metal2 -1642 -357 -1642 -357 1 clk
rlabel polycontact -1592 15 -1592 15 1 Y0
rlabel polycontact -1594 -141 -1594 -141 1 Y1
rlabel polycontact -1594 -349 -1594 -349 1 X0
rlabel polycontact -1597 -572 -1597 -572 1 X1
rlabel metal2 -101 -225 -101 -225 1 S1
rlabel metal1 -104 -207 -104 -207 1 C1
rlabel metal1 291 -208 291 -208 1 C2
rlabel metal2 -1361 15 -1361 15 1 Y0out
rlabel metal2 -1368 -141 -1368 -141 1 Y1out
rlabel metal2 -1368 -349 -1368 -349 1 X0out
rlabel metal2 -1372 -572 -1372 -572 1 X1out
rlabel metal2 326 -225 326 -225 1 S2
rlabel metal1 -78 -916 -78 -916 1 sum1
rlabel metal1 333 -931 333 -931 1 sum0
rlabel metal1 -941 -934 -941 -934 1 sum3
rlabel metal1 -552 -916 -552 -916 1 sum2
rlabel metal1 -1246 -661 -1246 -661 1 A1
rlabel polycontact -706 -661 -706 -661 1 Cin2
rlabel polycontact -790 -417 -790 -417 1 B
rlabel metal2 -494 -432 -494 -432 1 s3
rlabel metal1 -104 -424 -104 -424 1 c4
rlabel metal2 -85 -436 -85 -436 1 s4
rlabel metal1 -933 -658 -933 -658 1 c5
rlabel metal2 -926 -676 -926 -676 1 s5
rlabel metal1 -551 -657 -551 -657 1 c6
rlabel metal2 -547 -675 -547 -675 1 s6
rlabel metal1 -506 -422 -506 -422 1 c3
<< end >>
